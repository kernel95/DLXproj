----------------------------------------------------------------------------------
-- Create Date: 27.04.2021
-- Module Name: zero_comparator type 
-- Project Name: DLX
-- Version: 1.0
-- Additional Comments: type of conditions
----------------------------------------------------------------------------------

package comparator_type is 
    type TYPE_COMP is (ZERO, EQ, NEQ, GE, GT, LE, LT);
end comparator_type;
