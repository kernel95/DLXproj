
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_nwords64_isize32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_nwords64_isize32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity adder_genericu_nbit32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end adder_genericu_nbit32_DW01_add_0;

architecture SYN_rpl of adder_genericu_nbit32_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1002 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1002, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity adder_generic_nbit32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end adder_generic_nbit32_DW01_add_0;

architecture SYN_rpl of adder_generic_nbit32_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1005 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1005, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32_DW01_add_4 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end window_rf_M4_N4_F4_NBIT32_DW01_add_4;

architecture SYN_rpl of window_rf_M4_N4_F4_NBIT32_DW01_add_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_4_port, SUM_5_port, SUM_31_port, SUM_30_port, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, n29, n30, n31, n32, n33, n34, n35, n36, n37, 
      n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52
      , n53, n54, n55, SUM_3_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, A(2), A(1), A(0) );
   
   U1 : XOR2_X1 port map( A => A(4), B => A(3), Z => SUM_4_port);
   U2 : XOR2_X1 port map( A => A(5), B => n30, Z => SUM_5_port);
   U3 : XNOR2_X1 port map( A => A(31), B => n55, ZN => SUM_31_port);
   U4 : XOR2_X1 port map( A => A(30), B => n54, Z => SUM_30_port);
   U5 : XOR2_X1 port map( A => A(6), B => n29, Z => SUM_6_port);
   U6 : XOR2_X1 port map( A => A(7), B => n31, Z => SUM_7_port);
   U7 : XOR2_X1 port map( A => A(8), B => n32, Z => SUM_8_port);
   U8 : XOR2_X1 port map( A => A(9), B => n33, Z => SUM_9_port);
   U9 : XOR2_X1 port map( A => A(10), B => n34, Z => SUM_10_port);
   U10 : XOR2_X1 port map( A => A(11), B => n35, Z => SUM_11_port);
   U11 : XOR2_X1 port map( A => A(12), B => n36, Z => SUM_12_port);
   U12 : XOR2_X1 port map( A => A(13), B => n37, Z => SUM_13_port);
   U13 : XOR2_X1 port map( A => A(14), B => n38, Z => SUM_14_port);
   U14 : XOR2_X1 port map( A => A(15), B => n39, Z => SUM_15_port);
   U15 : XOR2_X1 port map( A => A(16), B => n40, Z => SUM_16_port);
   U16 : XOR2_X1 port map( A => A(17), B => n41, Z => SUM_17_port);
   U17 : XOR2_X1 port map( A => A(18), B => n42, Z => SUM_18_port);
   U18 : XOR2_X1 port map( A => A(19), B => n43, Z => SUM_19_port);
   U19 : XOR2_X1 port map( A => A(20), B => n44, Z => SUM_20_port);
   U20 : XOR2_X1 port map( A => A(21), B => n45, Z => SUM_21_port);
   U21 : XOR2_X1 port map( A => A(22), B => n46, Z => SUM_22_port);
   U22 : XOR2_X1 port map( A => A(23), B => n47, Z => SUM_23_port);
   U23 : XOR2_X1 port map( A => A(24), B => n48, Z => SUM_24_port);
   U24 : XOR2_X1 port map( A => A(25), B => n49, Z => SUM_25_port);
   U25 : XOR2_X1 port map( A => A(26), B => n50, Z => SUM_26_port);
   U26 : XOR2_X1 port map( A => A(27), B => n51, Z => SUM_27_port);
   U27 : XOR2_X1 port map( A => A(28), B => n52, Z => SUM_28_port);
   U28 : XOR2_X1 port map( A => A(29), B => n53, Z => SUM_29_port);
   U29 : NAND2_X1 port map( A1 => A(30), A2 => n54, ZN => n55);
   U30 : AND2_X1 port map( A1 => A(5), A2 => n30, ZN => n29);
   U31 : AND2_X1 port map( A1 => A(4), A2 => A(3), ZN => n30);
   U32 : AND2_X1 port map( A1 => A(6), A2 => n29, ZN => n31);
   U33 : AND2_X1 port map( A1 => A(7), A2 => n31, ZN => n32);
   U34 : AND2_X1 port map( A1 => A(8), A2 => n32, ZN => n33);
   U35 : AND2_X1 port map( A1 => A(9), A2 => n33, ZN => n34);
   U36 : AND2_X1 port map( A1 => A(10), A2 => n34, ZN => n35);
   U37 : AND2_X1 port map( A1 => A(11), A2 => n35, ZN => n36);
   U38 : AND2_X1 port map( A1 => A(12), A2 => n36, ZN => n37);
   U39 : AND2_X1 port map( A1 => A(13), A2 => n37, ZN => n38);
   U40 : AND2_X1 port map( A1 => A(14), A2 => n38, ZN => n39);
   U41 : AND2_X1 port map( A1 => A(15), A2 => n39, ZN => n40);
   U42 : AND2_X1 port map( A1 => A(16), A2 => n40, ZN => n41);
   U43 : AND2_X1 port map( A1 => A(17), A2 => n41, ZN => n42);
   U44 : AND2_X1 port map( A1 => A(18), A2 => n42, ZN => n43);
   U45 : AND2_X1 port map( A1 => A(19), A2 => n43, ZN => n44);
   U46 : AND2_X1 port map( A1 => A(20), A2 => n44, ZN => n45);
   U47 : AND2_X1 port map( A1 => A(21), A2 => n45, ZN => n46);
   U48 : AND2_X1 port map( A1 => A(22), A2 => n46, ZN => n47);
   U49 : AND2_X1 port map( A1 => A(23), A2 => n47, ZN => n48);
   U50 : AND2_X1 port map( A1 => A(24), A2 => n48, ZN => n49);
   U51 : AND2_X1 port map( A1 => A(25), A2 => n49, ZN => n50);
   U52 : AND2_X1 port map( A1 => A(26), A2 => n50, ZN => n51);
   U53 : AND2_X1 port map( A1 => A(27), A2 => n51, ZN => n52);
   U54 : AND2_X1 port map( A1 => A(28), A2 => n52, ZN => n53);
   U55 : AND2_X1 port map( A1 => A(29), A2 => n53, ZN => n54);
   U56 : INV_X1 port map( A => A(3), ZN => SUM_3_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32_DW01_sub_4 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end window_rf_M4_N4_F4_NBIT32_DW01_sub_4;

architecture SYN_rpl of window_rf_M4_N4_F4_NBIT32_DW01_sub_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, carry_31_port, carry_30_port, 
      carry_29_port, carry_28_port, carry_27_port, carry_26_port, carry_25_port
      , carry_24_port, carry_23_port, carry_22_port, carry_21_port, 
      carry_20_port, carry_19_port, carry_18_port, carry_17_port, carry_16_port
      , carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, n1, n2, n3, DIFF_3_port, n_1074 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, n_1074, 
      A(1), A(0) );
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => carry_6_port);
   U2 : INV_X1 port map( A => carry_5_port, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n1, A2 => DIFF_3_port, ZN => carry_5_port);
   U4 : INV_X1 port map( A => A(3), ZN => DIFF_3_port);
   U5 : XNOR2_X1 port map( A => A(4), B => A(3), ZN => DIFF_4_port);
   U6 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U7 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port);
   U8 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port);
   U9 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port);
   U10 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U11 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U12 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U13 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U14 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U15 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U16 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U17 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port)
                           ;
   U19 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port)
                           ;
   U20 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port)
                           ;
   U21 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port)
                           ;
   U22 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port)
                           ;
   U23 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port)
                           ;
   U24 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port)
                           ;
   U25 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port)
                           ;
   U26 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port)
                           ;
   U27 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port)
                           ;
   U28 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U29 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U30 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U31 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U32 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port)
                           ;
   U33 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U34 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U35 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U36 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U37 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U38 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U39 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U40 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U41 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U42 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U43 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U44 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U45 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U46 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U47 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U48 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U49 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U50 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U51 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U52 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U53 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U54 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U55 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U56 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U57 : OR2_X1 port map( A1 => A(30), A2 => carry_30_port, ZN => carry_31_port
                           );
   U58 : INV_X1 port map( A => A(4), ZN => n1);
   U59 : INV_X1 port map( A => A(5), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32_DW01_sub_3 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end window_rf_M4_N4_F4_NBIT32_DW01_sub_3;

architecture SYN_rpl of window_rf_M4_N4_F4_NBIT32_DW01_sub_3 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, carry_31_port, carry_30_port, 
      carry_29_port, carry_28_port, carry_27_port, carry_26_port, carry_25_port
      , carry_24_port, carry_23_port, carry_22_port, carry_21_port, 
      carry_20_port, carry_19_port, carry_18_port, carry_17_port, carry_16_port
      , carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, DIFF_3_port : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, A(2), 
      A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U2 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U3 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U4 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U5 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U6 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port);
   U7 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port);
   U8 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port);
   U9 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port);
   U10 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port)
                           ;
   U11 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port)
                           ;
   U12 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port)
                           ;
   U13 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port)
                           ;
   U14 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port)
                           ;
   U15 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port)
                           ;
   U16 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U17 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U19 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U20 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U21 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U22 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U23 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U24 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port)
                           ;
   U25 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port)
                           ;
   U26 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port)
                           ;
   U27 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port)
                           ;
   U28 : XNOR2_X1 port map( A => A(4), B => A(3), ZN => DIFF_4_port);
   U29 : INV_X1 port map( A => A(3), ZN => DIFF_3_port);
   U30 : OR2_X1 port map( A1 => A(4), A2 => A(3), ZN => carry_5_port);
   U31 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U32 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U33 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U34 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U35 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U36 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U37 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U38 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U39 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U40 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U41 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U42 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U43 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U44 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U45 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U46 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U47 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U48 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U49 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U50 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U51 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U52 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U53 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U54 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U55 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U56 : OR2_X1 port map( A1 => A(30), A2 => carry_30_port, ZN => carry_31_port
                           );

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32_DW01_add_3 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end window_rf_M4_N4_F4_NBIT32_DW01_add_3;

architecture SYN_rpl of window_rf_M4_N4_F4_NBIT32_DW01_add_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, n3 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n3, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM(5));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U3 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n3);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32_DW01_add_2 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end window_rf_M4_N4_F4_NBIT32_DW01_add_2;

architecture SYN_rpl of window_rf_M4_N4_F4_NBIT32_DW01_add_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, n3 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n3, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM(5));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U3 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n3);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32_DW01_add_1 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end window_rf_M4_N4_F4_NBIT32_DW01_add_1;

architecture SYN_rpl of window_rf_M4_N4_F4_NBIT32_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, n3 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n3, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM(5));
   U3 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n3);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end window_rf_M4_N4_F4_NBIT32_DW01_add_0;

architecture SYN_rpl of window_rf_M4_N4_F4_NBIT32_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_4_port, SUM_5_port, SUM_31_port, SUM_30_port, SUM_6_port, 
      SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, SUM_25_port, 
      SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, 
      SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, 
      SUM_14_port, SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, 
      SUM_9_port, SUM_8_port, SUM_7_port, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, SUM_3_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, A(2), A(1), A(0) );
   
   U1 : XOR2_X1 port map( A => A(4), B => A(3), Z => SUM_4_port);
   U2 : XOR2_X1 port map( A => A(5), B => n30, Z => SUM_5_port);
   U3 : XNOR2_X1 port map( A => A(31), B => n55, ZN => SUM_31_port);
   U4 : XOR2_X1 port map( A => A(30), B => n54, Z => SUM_30_port);
   U5 : XOR2_X1 port map( A => A(6), B => n29, Z => SUM_6_port);
   U6 : XOR2_X1 port map( A => A(29), B => n53, Z => SUM_29_port);
   U7 : XOR2_X1 port map( A => A(28), B => n52, Z => SUM_28_port);
   U8 : XOR2_X1 port map( A => A(27), B => n51, Z => SUM_27_port);
   U9 : XOR2_X1 port map( A => A(26), B => n50, Z => SUM_26_port);
   U10 : XOR2_X1 port map( A => A(25), B => n49, Z => SUM_25_port);
   U11 : XOR2_X1 port map( A => A(24), B => n48, Z => SUM_24_port);
   U12 : XOR2_X1 port map( A => A(23), B => n47, Z => SUM_23_port);
   U13 : XOR2_X1 port map( A => A(22), B => n46, Z => SUM_22_port);
   U14 : XOR2_X1 port map( A => A(21), B => n45, Z => SUM_21_port);
   U15 : XOR2_X1 port map( A => A(20), B => n44, Z => SUM_20_port);
   U16 : XOR2_X1 port map( A => A(19), B => n43, Z => SUM_19_port);
   U17 : XOR2_X1 port map( A => A(18), B => n42, Z => SUM_18_port);
   U18 : XOR2_X1 port map( A => A(17), B => n41, Z => SUM_17_port);
   U19 : XOR2_X1 port map( A => A(16), B => n40, Z => SUM_16_port);
   U20 : XOR2_X1 port map( A => A(15), B => n39, Z => SUM_15_port);
   U21 : XOR2_X1 port map( A => A(14), B => n38, Z => SUM_14_port);
   U22 : XOR2_X1 port map( A => A(13), B => n37, Z => SUM_13_port);
   U23 : XOR2_X1 port map( A => A(12), B => n36, Z => SUM_12_port);
   U24 : XOR2_X1 port map( A => A(11), B => n35, Z => SUM_11_port);
   U25 : XOR2_X1 port map( A => A(10), B => n34, Z => SUM_10_port);
   U26 : XOR2_X1 port map( A => A(9), B => n33, Z => SUM_9_port);
   U27 : XOR2_X1 port map( A => A(8), B => n32, Z => SUM_8_port);
   U28 : XOR2_X1 port map( A => A(7), B => n31, Z => SUM_7_port);
   U29 : AND2_X1 port map( A1 => A(5), A2 => n30, ZN => n29);
   U30 : AND2_X1 port map( A1 => A(4), A2 => A(3), ZN => n30);
   U31 : NAND2_X1 port map( A1 => A(30), A2 => n54, ZN => n55);
   U32 : INV_X1 port map( A => A(3), ZN => SUM_3_port);
   U33 : AND2_X1 port map( A1 => A(6), A2 => n29, ZN => n31);
   U34 : AND2_X1 port map( A1 => A(7), A2 => n31, ZN => n32);
   U35 : AND2_X1 port map( A1 => A(8), A2 => n32, ZN => n33);
   U36 : AND2_X1 port map( A1 => A(9), A2 => n33, ZN => n34);
   U37 : AND2_X1 port map( A1 => A(10), A2 => n34, ZN => n35);
   U38 : AND2_X1 port map( A1 => A(11), A2 => n35, ZN => n36);
   U39 : AND2_X1 port map( A1 => A(12), A2 => n36, ZN => n37);
   U40 : AND2_X1 port map( A1 => A(13), A2 => n37, ZN => n38);
   U41 : AND2_X1 port map( A1 => A(14), A2 => n38, ZN => n39);
   U42 : AND2_X1 port map( A1 => A(15), A2 => n39, ZN => n40);
   U43 : AND2_X1 port map( A1 => A(16), A2 => n40, ZN => n41);
   U44 : AND2_X1 port map( A1 => A(17), A2 => n41, ZN => n42);
   U45 : AND2_X1 port map( A1 => A(18), A2 => n42, ZN => n43);
   U46 : AND2_X1 port map( A1 => A(19), A2 => n43, ZN => n44);
   U47 : AND2_X1 port map( A1 => A(20), A2 => n44, ZN => n45);
   U48 : AND2_X1 port map( A1 => A(21), A2 => n45, ZN => n46);
   U49 : AND2_X1 port map( A1 => A(22), A2 => n46, ZN => n47);
   U50 : AND2_X1 port map( A1 => A(23), A2 => n47, ZN => n48);
   U51 : AND2_X1 port map( A1 => A(24), A2 => n48, ZN => n49);
   U52 : AND2_X1 port map( A1 => A(25), A2 => n49, ZN => n50);
   U53 : AND2_X1 port map( A1 => A(26), A2 => n50, ZN => n51);
   U54 : AND2_X1 port map( A1 => A(27), A2 => n51, ZN => n52);
   U55 : AND2_X1 port map( A1 => A(28), A2 => n52, ZN => n53);
   U56 : AND2_X1 port map( A1 => A(29), A2 => n53, ZN => n54);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity comparator_addr_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_addr_DW01_cmp6_0;

architecture SYN_rpl of comparator_addr_DW01_cmp6_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A(1), ZN => n2);
   U2 : INV_X1 port map( A => A(0), ZN => n3);
   U3 : INV_X1 port map( A => B(1), ZN => n1);
   U4 : NOR4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => EQ);
   U5 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n7);
   U6 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n11);
   U7 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n10);
   U8 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n9);
   U9 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n8);
   U10 : NAND4_X1 port map( A1 => n12, A2 => n13, A3 => n14, A4 => n15, ZN => 
                           n6);
   U11 : OAI22_X1 port map( A1 => n16, A2 => n2, B1 => B(1), B2 => n16, ZN => 
                           n15);
   U12 : AND2_X1 port map( A1 => B(0), A2 => n3, ZN => n16);
   U13 : OAI22_X1 port map( A1 => A(1), A2 => n17, B1 => n17, B2 => n1, ZN => 
                           n14);
   U14 : NOR2_X1 port map( A1 => n3, A2 => B(0), ZN => n17);
   U15 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n13);
   U16 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n12);
   U17 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n5);
   U18 : NOR4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => 
                           n19);
   U19 : XOR2_X1 port map( A => B(10), B => A(10), Z => n23);
   U20 : XOR2_X1 port map( A => B(9), B => A(9), Z => n22);
   U21 : XOR2_X1 port map( A => B(8), B => A(8), Z => n21);
   U22 : XOR2_X1 port map( A => B(7), B => A(7), Z => n20);
   U23 : NOR4_X1 port map( A1 => n24, A2 => n25, A3 => n26, A4 => n27, ZN => 
                           n18);
   U24 : XOR2_X1 port map( A => B(14), B => A(14), Z => n27);
   U25 : XOR2_X1 port map( A => B(13), B => A(13), Z => n26);
   U26 : XOR2_X1 port map( A => B(12), B => A(12), Z => n25);
   U27 : XOR2_X1 port map( A => B(11), B => A(11), Z => n24);
   U28 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n4);
   U29 : NOR4_X1 port map( A1 => n32, A2 => n33, A3 => n34, A4 => n35, ZN => 
                           n31);
   U30 : XOR2_X1 port map( A => B(18), B => A(18), Z => n35);
   U31 : XOR2_X1 port map( A => B(17), B => A(17), Z => n34);
   U32 : XOR2_X1 port map( A => B(16), B => A(16), Z => n33);
   U33 : XOR2_X1 port map( A => B(15), B => A(15), Z => n32);
   U34 : NOR4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => 
                           n30);
   U35 : XOR2_X1 port map( A => B(22), B => A(22), Z => n39);
   U36 : XOR2_X1 port map( A => B(21), B => A(21), Z => n38);
   U37 : XOR2_X1 port map( A => B(20), B => A(20), Z => n37);
   U38 : XOR2_X1 port map( A => B(19), B => A(19), Z => n36);
   U39 : NOR4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n29);
   U40 : XOR2_X1 port map( A => B(26), B => A(26), Z => n43);
   U41 : XOR2_X1 port map( A => B(25), B => A(25), Z => n42);
   U42 : XOR2_X1 port map( A => B(24), B => A(24), Z => n41);
   U43 : XOR2_X1 port map( A => B(23), B => A(23), Z => n40);
   U44 : NOR4_X1 port map( A1 => n44, A2 => n45, A3 => n46, A4 => n47, ZN => 
                           n28);
   U45 : XOR2_X1 port map( A => B(30), B => A(30), Z => n47);
   U46 : XOR2_X1 port map( A => B(29), B => A(29), Z => n46);
   U47 : XOR2_X1 port map( A => B(28), B => A(28), Z => n45);
   U48 : XOR2_X1 port map( A => B(27), B => A(27), Z => n44);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity zero_comparator_N32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end zero_comparator_N32_DW01_cmp6_0;

architecture SYN_rpl of zero_comparator_N32_DW01_cmp6_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GT_port, n202, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201 : std_logic;

begin
   GT <= GT_port;
   
   U1 : INV_X1 port map( A => n141, ZN => n29);
   U2 : INV_X1 port map( A => n129, ZN => n25);
   U3 : INV_X1 port map( A => n117, ZN => n21);
   U4 : INV_X1 port map( A => n105, ZN => n17);
   U5 : INV_X1 port map( A => n93, ZN => n13);
   U6 : INV_X1 port map( A => n81, ZN => n9);
   U7 : INV_X1 port map( A => n126, ZN => n24);
   U8 : INV_X1 port map( A => n114, ZN => n20);
   U9 : INV_X1 port map( A => n102, ZN => n16);
   U10 : INV_X1 port map( A => n90, ZN => n12);
   U11 : INV_X1 port map( A => n78, ZN => n8);
   U12 : INV_X1 port map( A => n143, ZN => n31);
   U13 : INV_X1 port map( A => n131, ZN => n27);
   U14 : INV_X1 port map( A => n119, ZN => n23);
   U15 : INV_X1 port map( A => n153, ZN => n33);
   U16 : INV_X1 port map( A => n140, ZN => n30);
   U17 : INV_X1 port map( A => n128, ZN => n26);
   U18 : INV_X1 port map( A => n116, ZN => n22);
   U19 : INV_X1 port map( A => n107, ZN => n19);
   U20 : INV_X1 port map( A => n95, ZN => n15);
   U21 : INV_X1 port map( A => n83, ZN => n11);
   U22 : INV_X1 port map( A => n104, ZN => n18);
   U23 : INV_X1 port map( A => n92, ZN => n14);
   U24 : INV_X1 port map( A => n80, ZN => n10);
   U25 : INV_X1 port map( A => n138, ZN => n28);
   U26 : INV_X1 port map( A => GT_port, ZN => n2);
   U27 : INV_X1 port map( A => B(1), ZN => n35);
   U28 : INV_X1 port map( A => B(30), ZN => n6);
   U29 : INV_X1 port map( A => n202, ZN => LT);
   U30 : INV_X1 port map( A => B(31), ZN => n4);
   U31 : INV_X1 port map( A => A(0), ZN => n64);
   U32 : INV_X1 port map( A => n67, ZN => n5);
   U33 : INV_X1 port map( A => A(30), ZN => n36);
   U34 : INV_X1 port map( A => n71, ZN => n7);
   U35 : INV_X1 port map( A => A(5), ZN => n60);
   U36 : INV_X1 port map( A => A(9), ZN => n56);
   U37 : INV_X1 port map( A => A(11), ZN => n54);
   U38 : INV_X1 port map( A => A(3), ZN => n62);
   U39 : INV_X1 port map( A => A(7), ZN => n58);
   U40 : INV_X1 port map( A => A(13), ZN => n52);
   U41 : INV_X1 port map( A => A(12), ZN => n53);
   U42 : INV_X1 port map( A => A(4), ZN => n61);
   U43 : INV_X1 port map( A => A(8), ZN => n57);
   U44 : INV_X1 port map( A => A(2), ZN => n63);
   U45 : INV_X1 port map( A => A(10), ZN => n55);
   U46 : INV_X1 port map( A => A(14), ZN => n51);
   U47 : INV_X1 port map( A => A(6), ZN => n59);
   U48 : INV_X1 port map( A => A(27), ZN => n39);
   U49 : INV_X1 port map( A => A(23), ZN => n43);
   U50 : INV_X1 port map( A => A(19), ZN => n47);
   U51 : INV_X1 port map( A => A(25), ZN => n41);
   U52 : INV_X1 port map( A => A(29), ZN => n37);
   U53 : INV_X1 port map( A => A(21), ZN => n45);
   U54 : INV_X1 port map( A => A(17), ZN => n49);
   U55 : INV_X1 port map( A => A(16), ZN => n50);
   U56 : INV_X1 port map( A => A(24), ZN => n42);
   U57 : INV_X1 port map( A => A(28), ZN => n38);
   U58 : INV_X1 port map( A => A(20), ZN => n46);
   U59 : INV_X1 port map( A => A(26), ZN => n40);
   U60 : INV_X1 port map( A => A(22), ZN => n44);
   U61 : INV_X1 port map( A => A(18), ZN => n48);
   U62 : INV_X1 port map( A => n201, ZN => n34);
   U63 : INV_X1 port map( A => n150, ZN => n32);
   U64 : INV_X1 port map( A => A(15), ZN => n1);
   U65 : NAND2_X1 port map( A1 => n2, A2 => n202, ZN => NE);
   U66 : AOI21_X1 port map( B1 => n65, B2 => n5, A => n66, ZN => n202);
   U67 : AOI22_X1 port map( A1 => B(30), A2 => n36, B1 => n68, B2 => n69, ZN =>
                           n67);
   U68 : AOI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n68);
   U69 : AOI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n70);
   U70 : AOI21_X1 port map( B1 => n76, B2 => n77, A => n78, ZN => n73);
   U71 : AOI21_X1 port map( B1 => n79, B2 => n9, A => n10, ZN => n76);
   U72 : AOI21_X1 port map( B1 => n82, B2 => n83, A => n84, ZN => n79);
   U73 : AOI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n82);
   U74 : AOI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n85);
   U75 : AOI21_X1 port map( B1 => n91, B2 => n13, A => n14, ZN => n88);
   U76 : AOI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n91);
   U77 : AOI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n94);
   U78 : AOI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => n97);
   U79 : AOI21_X1 port map( B1 => n103, B2 => n17, A => n18, ZN => n100);
   U80 : AOI21_X1 port map( B1 => n106, B2 => n107, A => n108, ZN => n103);
   U81 : AOI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n106);
   U82 : AOI21_X1 port map( B1 => n112, B2 => n113, A => n114, ZN => n109);
   U83 : AOI21_X1 port map( B1 => n115, B2 => n21, A => n22, ZN => n112);
   U84 : AOI21_X1 port map( B1 => n118, B2 => n119, A => n120, ZN => n115);
   U85 : AOI21_X1 port map( B1 => n121, B2 => n122, A => n123, ZN => n118);
   U86 : AOI21_X1 port map( B1 => n124, B2 => n125, A => n126, ZN => n121);
   U87 : AOI21_X1 port map( B1 => n127, B2 => n25, A => n26, ZN => n124);
   U88 : AOI21_X1 port map( B1 => n130, B2 => n131, A => n132, ZN => n127);
   U89 : AOI21_X1 port map( B1 => n133, B2 => n134, A => n135, ZN => n130);
   U90 : AOI21_X1 port map( B1 => n136, B2 => n137, A => n138, ZN => n133);
   U91 : AOI21_X1 port map( B1 => n139, B2 => n29, A => n30, ZN => n136);
   U92 : AOI21_X1 port map( B1 => n142, B2 => n143, A => n144, ZN => n139);
   U93 : AOI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n142);
   U94 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n145);
   U95 : AOI21_X1 port map( B1 => n151, B2 => n152, A => n33, ZN => n148);
   U96 : AOI22_X1 port map( A1 => n154, A2 => n35, B1 => A(1), B2 => n155, ZN 
                           => n151);
   U97 : OR2_X1 port map( A1 => n155, A2 => A(1), ZN => n154);
   U98 : NAND2_X1 port map( A1 => B(0), A2 => n64, ZN => n155);
   U99 : OAI21_X1 port map( B1 => n66, B2 => n156, A => n65, ZN => GT_port);
   U100 : NAND2_X1 port map( A1 => A(31), A2 => n4, ZN => n65);
   U101 : AOI22_X1 port map( A1 => A(30), A2 => n6, B1 => n157, B2 => n69, ZN 
                           => n156);
   U102 : XOR2_X1 port map( A => A(30), B => n6, Z => n69);
   U103 : AOI21_X1 port map( B1 => n158, B2 => n159, A => n7, ZN => n157);
   U104 : NAND2_X1 port map( A1 => B(29), A2 => n37, ZN => n71);
   U105 : OAI211_X1 port map( C1 => n160, C2 => n161, A => n77, B => n74, ZN =>
                           n159);
   U106 : NOR2_X1 port map( A1 => n162, A2 => n75, ZN => n74);
   U107 : AND2_X1 port map( A1 => B(28), A2 => n38, ZN => n75);
   U108 : NAND2_X1 port map( A1 => B(27), A2 => n39, ZN => n77);
   U109 : NAND2_X1 port map( A1 => n8, A2 => n163, ZN => n161);
   U110 : NOR2_X1 port map( A1 => n39, A2 => B(27), ZN => n78);
   U111 : AOI211_X1 port map( C1 => n164, C2 => n165, A => n81, B => n11, ZN =>
                           n160);
   U112 : NAND2_X1 port map( A1 => B(25), A2 => n41, ZN => n83);
   U113 : NAND2_X1 port map( A1 => n163, A2 => n80, ZN => n81);
   U114 : NAND2_X1 port map( A1 => B(26), A2 => n40, ZN => n80);
   U115 : OR2_X1 port map( A1 => n40, A2 => B(26), ZN => n163);
   U116 : OAI211_X1 port map( C1 => n166, C2 => n167, A => n89, B => n86, ZN =>
                           n165);
   U117 : NOR2_X1 port map( A1 => n168, A2 => n87, ZN => n86);
   U118 : AND2_X1 port map( A1 => B(24), A2 => n42, ZN => n87);
   U119 : NAND2_X1 port map( A1 => B(23), A2 => n43, ZN => n89);
   U120 : NAND2_X1 port map( A1 => n12, A2 => n169, ZN => n167);
   U121 : NOR2_X1 port map( A1 => n43, A2 => B(23), ZN => n90);
   U122 : AOI211_X1 port map( C1 => n170, C2 => n171, A => n93, B => n15, ZN =>
                           n166);
   U123 : NAND2_X1 port map( A1 => B(21), A2 => n45, ZN => n95);
   U124 : NAND2_X1 port map( A1 => n169, A2 => n92, ZN => n93);
   U125 : NAND2_X1 port map( A1 => B(22), A2 => n44, ZN => n92);
   U126 : OR2_X1 port map( A1 => n44, A2 => B(22), ZN => n169);
   U127 : OAI211_X1 port map( C1 => n172, C2 => n173, A => n101, B => n98, ZN 
                           => n171);
   U128 : NOR2_X1 port map( A1 => n174, A2 => n99, ZN => n98);
   U129 : AND2_X1 port map( A1 => B(20), A2 => n46, ZN => n99);
   U130 : NAND2_X1 port map( A1 => B(19), A2 => n47, ZN => n101);
   U131 : NAND2_X1 port map( A1 => n16, A2 => n175, ZN => n173);
   U132 : NOR2_X1 port map( A1 => n47, A2 => B(19), ZN => n102);
   U133 : AOI211_X1 port map( C1 => n176, C2 => n177, A => n105, B => n19, ZN 
                           => n172);
   U134 : NAND2_X1 port map( A1 => B(17), A2 => n49, ZN => n107);
   U135 : NAND2_X1 port map( A1 => n175, A2 => n104, ZN => n105);
   U136 : NAND2_X1 port map( A1 => B(18), A2 => n48, ZN => n104);
   U137 : OR2_X1 port map( A1 => n48, A2 => B(18), ZN => n175);
   U138 : OAI211_X1 port map( C1 => n178, C2 => n179, A => n113, B => n110, ZN 
                           => n177);
   U139 : NOR2_X1 port map( A1 => n180, A2 => n111, ZN => n110);
   U140 : AND2_X1 port map( A1 => B(16), A2 => n50, ZN => n111);
   U141 : NAND2_X1 port map( A1 => B(15), A2 => n1, ZN => n113);
   U142 : NAND2_X1 port map( A1 => n20, A2 => n181, ZN => n179);
   U143 : NOR2_X1 port map( A1 => n1, A2 => B(15), ZN => n114);
   U144 : AOI211_X1 port map( C1 => n182, C2 => n183, A => n117, B => n23, ZN 
                           => n178);
   U145 : NAND2_X1 port map( A1 => B(13), A2 => n52, ZN => n119);
   U146 : NAND2_X1 port map( A1 => n181, A2 => n116, ZN => n117);
   U147 : NAND2_X1 port map( A1 => B(14), A2 => n51, ZN => n116);
   U148 : OR2_X1 port map( A1 => n51, A2 => B(14), ZN => n181);
   U149 : OAI211_X1 port map( C1 => n184, C2 => n185, A => n125, B => n122, ZN 
                           => n183);
   U150 : NOR2_X1 port map( A1 => n186, A2 => n123, ZN => n122);
   U151 : AND2_X1 port map( A1 => B(12), A2 => n53, ZN => n123);
   U152 : NAND2_X1 port map( A1 => B(11), A2 => n54, ZN => n125);
   U153 : NAND2_X1 port map( A1 => n24, A2 => n187, ZN => n185);
   U154 : NOR2_X1 port map( A1 => n54, A2 => B(11), ZN => n126);
   U155 : AOI211_X1 port map( C1 => n188, C2 => n189, A => n129, B => n27, ZN 
                           => n184);
   U156 : NAND2_X1 port map( A1 => B(9), A2 => n56, ZN => n131);
   U157 : NAND2_X1 port map( A1 => n187, A2 => n128, ZN => n129);
   U158 : NAND2_X1 port map( A1 => B(10), A2 => n55, ZN => n128);
   U159 : OR2_X1 port map( A1 => n55, A2 => B(10), ZN => n187);
   U160 : OAI211_X1 port map( C1 => n190, C2 => n191, A => n137, B => n134, ZN 
                           => n189);
   U161 : NOR2_X1 port map( A1 => n192, A2 => n135, ZN => n134);
   U162 : AND2_X1 port map( A1 => B(8), A2 => n57, ZN => n135);
   U163 : NAND2_X1 port map( A1 => B(7), A2 => n58, ZN => n137);
   U164 : NAND2_X1 port map( A1 => n28, A2 => n193, ZN => n191);
   U165 : NOR2_X1 port map( A1 => n58, A2 => B(7), ZN => n138);
   U166 : AOI211_X1 port map( C1 => n194, C2 => n195, A => n141, B => n31, ZN 
                           => n190);
   U167 : NAND2_X1 port map( A1 => B(5), A2 => n60, ZN => n143);
   U168 : NAND2_X1 port map( A1 => n193, A2 => n140, ZN => n141);
   U169 : NAND2_X1 port map( A1 => B(6), A2 => n59, ZN => n140);
   U170 : OR2_X1 port map( A1 => n59, A2 => B(6), ZN => n193);
   U171 : NAND3_X1 port map( A1 => n196, A2 => n149, A3 => n146, ZN => n195);
   U172 : NOR2_X1 port map( A1 => n197, A2 => n147, ZN => n146);
   U173 : AND2_X1 port map( A1 => B(4), A2 => n61, ZN => n147);
   U174 : NAND2_X1 port map( A1 => B(3), A2 => n62, ZN => n149);
   U175 : NAND3_X1 port map( A1 => n32, A2 => n198, A3 => n199, ZN => n196);
   U176 : OAI211_X1 port map( C1 => A(1), C2 => n200, A => n34, B => n152, ZN 
                           => n199);
   U177 : AND2_X1 port map( A1 => n198, A2 => n153, ZN => n152);
   U178 : NAND2_X1 port map( A1 => B(2), A2 => n63, ZN => n153);
   U179 : AOI21_X1 port map( B1 => A(1), B2 => n200, A => n35, ZN => n201);
   U180 : NOR2_X1 port map( A1 => n64, A2 => B(0), ZN => n200);
   U181 : OR2_X1 port map( A1 => n63, A2 => B(2), ZN => n198);
   U182 : NOR2_X1 port map( A1 => n62, A2 => B(3), ZN => n150);
   U183 : NOR2_X1 port map( A1 => n197, A2 => n144, ZN => n194);
   U184 : NOR2_X1 port map( A1 => n60, A2 => B(5), ZN => n144);
   U185 : NOR2_X1 port map( A1 => n61, A2 => B(4), ZN => n197);
   U186 : NOR2_X1 port map( A1 => n192, A2 => n132, ZN => n188);
   U187 : NOR2_X1 port map( A1 => n56, A2 => B(9), ZN => n132);
   U188 : NOR2_X1 port map( A1 => n57, A2 => B(8), ZN => n192);
   U189 : NOR2_X1 port map( A1 => n186, A2 => n120, ZN => n182);
   U190 : NOR2_X1 port map( A1 => n52, A2 => B(13), ZN => n120);
   U191 : NOR2_X1 port map( A1 => n53, A2 => B(12), ZN => n186);
   U192 : NOR2_X1 port map( A1 => n180, A2 => n108, ZN => n176);
   U193 : NOR2_X1 port map( A1 => n49, A2 => B(17), ZN => n108);
   U194 : NOR2_X1 port map( A1 => n50, A2 => B(16), ZN => n180);
   U195 : NOR2_X1 port map( A1 => n174, A2 => n96, ZN => n170);
   U196 : NOR2_X1 port map( A1 => n45, A2 => B(21), ZN => n96);
   U197 : NOR2_X1 port map( A1 => n46, A2 => B(20), ZN => n174);
   U198 : NOR2_X1 port map( A1 => n168, A2 => n84, ZN => n164);
   U199 : NOR2_X1 port map( A1 => n41, A2 => B(25), ZN => n84);
   U200 : NOR2_X1 port map( A1 => n42, A2 => B(24), ZN => n168);
   U201 : NOR2_X1 port map( A1 => n162, A2 => n72, ZN => n158);
   U202 : NOR2_X1 port map( A1 => n37, A2 => B(29), ZN => n72);
   U203 : NOR2_X1 port map( A1 => n38, A2 => B(28), ZN => n162);
   U204 : NOR2_X1 port map( A1 => n4, A2 => A(31), ZN => n66);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_216 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_216;

architecture SYN_Behavioral of or2_216 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_215 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_215;

architecture SYN_Behavioral of or2_215 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_214 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_214;

architecture SYN_Behavioral of or2_214 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_213 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_213;

architecture SYN_Behavioral of or2_213 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_212 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_212;

architecture SYN_Behavioral of or2_212 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_211 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_211;

architecture SYN_Behavioral of or2_211 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_210 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_210;

architecture SYN_Behavioral of or2_210 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_209 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_209;

architecture SYN_Behavioral of or2_209 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_208 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_208;

architecture SYN_Behavioral of or2_208 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_207 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_207;

architecture SYN_Behavioral of or2_207 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_206 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_206;

architecture SYN_Behavioral of or2_206 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_205 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_205;

architecture SYN_Behavioral of or2_205 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_204 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_204;

architecture SYN_Behavioral of or2_204 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_203 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_203;

architecture SYN_Behavioral of or2_203 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_202 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_202;

architecture SYN_Behavioral of or2_202 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_201 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_201;

architecture SYN_Behavioral of or2_201 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_200 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_200;

architecture SYN_Behavioral of or2_200 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_199 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_199;

architecture SYN_Behavioral of or2_199 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_198 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_198;

architecture SYN_Behavioral of or2_198 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_197 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_197;

architecture SYN_Behavioral of or2_197 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_196 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_196;

architecture SYN_Behavioral of or2_196 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_195 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_195;

architecture SYN_Behavioral of or2_195 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_194 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_194;

architecture SYN_Behavioral of or2_194 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_193 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_193;

architecture SYN_Behavioral of or2_193 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_192 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_192;

architecture SYN_Behavioral of or2_192 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_191 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_191;

architecture SYN_Behavioral of or2_191 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_190 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_190;

architecture SYN_Behavioral of or2_190 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_189 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_189;

architecture SYN_Behavioral of or2_189 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_188 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_188;

architecture SYN_Behavioral of or2_188 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_187 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_187;

architecture SYN_Behavioral of or2_187 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_186 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_186;

architecture SYN_Behavioral of or2_186 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_185 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_185;

architecture SYN_Behavioral of or2_185 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_184 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_184;

architecture SYN_Behavioral of or2_184 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_183 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_183;

architecture SYN_Behavioral of or2_183 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_182 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_182;

architecture SYN_Behavioral of or2_182 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_181 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_181;

architecture SYN_Behavioral of or2_181 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_180 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_180;

architecture SYN_Behavioral of or2_180 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_179 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_179;

architecture SYN_Behavioral of or2_179 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_178 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_178;

architecture SYN_Behavioral of or2_178 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_177 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_177;

architecture SYN_Behavioral of or2_177 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_176 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_176;

architecture SYN_Behavioral of or2_176 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_175 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_175;

architecture SYN_Behavioral of or2_175 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_174 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_174;

architecture SYN_Behavioral of or2_174 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_173 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_173;

architecture SYN_Behavioral of or2_173 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_172 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_172;

architecture SYN_Behavioral of or2_172 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_171 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_171;

architecture SYN_Behavioral of or2_171 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_170 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_170;

architecture SYN_Behavioral of or2_170 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_169 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_169;

architecture SYN_Behavioral of or2_169 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_168 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_168;

architecture SYN_Behavioral of or2_168 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_167 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_167;

architecture SYN_Behavioral of or2_167 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_166 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_166;

architecture SYN_Behavioral of or2_166 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_165 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_165;

architecture SYN_Behavioral of or2_165 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_164 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_164;

architecture SYN_Behavioral of or2_164 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_163 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_163;

architecture SYN_Behavioral of or2_163 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_162 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_162;

architecture SYN_Behavioral of or2_162 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_161 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_161;

architecture SYN_Behavioral of or2_161 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_160 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_160;

architecture SYN_Behavioral of or2_160 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_159 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_159;

architecture SYN_Behavioral of or2_159 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_158 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_158;

architecture SYN_Behavioral of or2_158 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_157 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_157;

architecture SYN_Behavioral of or2_157 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_156 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_156;

architecture SYN_Behavioral of or2_156 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_155 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_155;

architecture SYN_Behavioral of or2_155 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_154 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_154;

architecture SYN_Behavioral of or2_154 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_153 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_153;

architecture SYN_Behavioral of or2_153 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_152 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_152;

architecture SYN_Behavioral of or2_152 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_151 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_151;

architecture SYN_Behavioral of or2_151 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_150 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_150;

architecture SYN_Behavioral of or2_150 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_149 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_149;

architecture SYN_Behavioral of or2_149 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_148 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_148;

architecture SYN_Behavioral of or2_148 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_147 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_147;

architecture SYN_Behavioral of or2_147 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_146 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_146;

architecture SYN_Behavioral of or2_146 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_145 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_145;

architecture SYN_Behavioral of or2_145 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_144 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_144;

architecture SYN_Behavioral of or2_144 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_143 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_143;

architecture SYN_Behavioral of or2_143 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_142 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_142;

architecture SYN_Behavioral of or2_142 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_141 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_141;

architecture SYN_Behavioral of or2_141 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_140 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_140;

architecture SYN_Behavioral of or2_140 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_139 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_139;

architecture SYN_Behavioral of or2_139 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_138 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_138;

architecture SYN_Behavioral of or2_138 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_137 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_137;

architecture SYN_Behavioral of or2_137 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_136 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_136;

architecture SYN_Behavioral of or2_136 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_135 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_135;

architecture SYN_Behavioral of or2_135 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_134 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_134;

architecture SYN_Behavioral of or2_134 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_133 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_133;

architecture SYN_Behavioral of or2_133 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_132 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_132;

architecture SYN_Behavioral of or2_132 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_131 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_131;

architecture SYN_Behavioral of or2_131 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_130 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_130;

architecture SYN_Behavioral of or2_130 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_129 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_129;

architecture SYN_Behavioral of or2_129 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_128 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_128;

architecture SYN_Behavioral of or2_128 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_127 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_127;

architecture SYN_Behavioral of or2_127 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_126 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_126;

architecture SYN_Behavioral of or2_126 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_125 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_125;

architecture SYN_Behavioral of or2_125 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_124 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_124;

architecture SYN_Behavioral of or2_124 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_123 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_123;

architecture SYN_Behavioral of or2_123 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_122 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_122;

architecture SYN_Behavioral of or2_122 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_121 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_121;

architecture SYN_Behavioral of or2_121 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_120 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_120;

architecture SYN_Behavioral of or2_120 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_119 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_119;

architecture SYN_Behavioral of or2_119 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_118 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_118;

architecture SYN_Behavioral of or2_118 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_117 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_117;

architecture SYN_Behavioral of or2_117 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_116 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_116;

architecture SYN_Behavioral of or2_116 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_115 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_115;

architecture SYN_Behavioral of or2_115 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_114 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_114;

architecture SYN_Behavioral of or2_114 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_113 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_113;

architecture SYN_Behavioral of or2_113 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_112 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_112;

architecture SYN_Behavioral of or2_112 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_111 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_111;

architecture SYN_Behavioral of or2_111 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_110 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_110;

architecture SYN_Behavioral of or2_110 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_109 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_109;

architecture SYN_Behavioral of or2_109 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_108 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_108;

architecture SYN_Behavioral of or2_108 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_107 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_107;

architecture SYN_Behavioral of or2_107 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_106 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_106;

architecture SYN_Behavioral of or2_106 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_105 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_105;

architecture SYN_Behavioral of or2_105 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_104 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_104;

architecture SYN_Behavioral of or2_104 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_103 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_103;

architecture SYN_Behavioral of or2_103 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_102 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_102;

architecture SYN_Behavioral of or2_102 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_101 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_101;

architecture SYN_Behavioral of or2_101 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_100 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_100;

architecture SYN_Behavioral of or2_100 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_99 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_99;

architecture SYN_Behavioral of or2_99 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_98 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_98;

architecture SYN_Behavioral of or2_98 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_97 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_97;

architecture SYN_Behavioral of or2_97 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_96 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_96;

architecture SYN_Behavioral of or2_96 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_95 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_95;

architecture SYN_Behavioral of or2_95 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_94 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_94;

architecture SYN_Behavioral of or2_94 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_93 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_93;

architecture SYN_Behavioral of or2_93 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_92 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_92;

architecture SYN_Behavioral of or2_92 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_91 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_91;

architecture SYN_Behavioral of or2_91 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_90 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_90;

architecture SYN_Behavioral of or2_90 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_89 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_89;

architecture SYN_Behavioral of or2_89 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_88 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_88;

architecture SYN_Behavioral of or2_88 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_87 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_87;

architecture SYN_Behavioral of or2_87 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_86 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_86;

architecture SYN_Behavioral of or2_86 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_85 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_85;

architecture SYN_Behavioral of or2_85 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_84 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_84;

architecture SYN_Behavioral of or2_84 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_83 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_83;

architecture SYN_Behavioral of or2_83 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_82 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_82;

architecture SYN_Behavioral of or2_82 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_81 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_81;

architecture SYN_Behavioral of or2_81 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_80 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_80;

architecture SYN_Behavioral of or2_80 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_79 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_79;

architecture SYN_Behavioral of or2_79 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_78 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_78;

architecture SYN_Behavioral of or2_78 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_77 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_77;

architecture SYN_Behavioral of or2_77 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_76 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_76;

architecture SYN_Behavioral of or2_76 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_75 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_75;

architecture SYN_Behavioral of or2_75 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_74 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_74;

architecture SYN_Behavioral of or2_74 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_73 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_73;

architecture SYN_Behavioral of or2_73 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_72 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_72;

architecture SYN_Behavioral of or2_72 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_71 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_71;

architecture SYN_Behavioral of or2_71 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_70 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_70;

architecture SYN_Behavioral of or2_70 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_69 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_69;

architecture SYN_Behavioral of or2_69 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_68 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_68;

architecture SYN_Behavioral of or2_68 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_67 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_67;

architecture SYN_Behavioral of or2_67 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_66 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_66;

architecture SYN_Behavioral of or2_66 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_65 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_65;

architecture SYN_Behavioral of or2_65 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_64 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_64;

architecture SYN_Behavioral of or2_64 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_63 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_63;

architecture SYN_Behavioral of or2_63 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_62 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_62;

architecture SYN_Behavioral of or2_62 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_61 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_61;

architecture SYN_Behavioral of or2_61 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_60 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_60;

architecture SYN_Behavioral of or2_60 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_59 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_59;

architecture SYN_Behavioral of or2_59 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_58 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_58;

architecture SYN_Behavioral of or2_58 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_57 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_57;

architecture SYN_Behavioral of or2_57 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_56 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_56;

architecture SYN_Behavioral of or2_56 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_55 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_55;

architecture SYN_Behavioral of or2_55 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_54 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_54;

architecture SYN_Behavioral of or2_54 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_53 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_53;

architecture SYN_Behavioral of or2_53 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_52 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_52;

architecture SYN_Behavioral of or2_52 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_51 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_51;

architecture SYN_Behavioral of or2_51 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_50 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_50;

architecture SYN_Behavioral of or2_50 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_49 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_49;

architecture SYN_Behavioral of or2_49 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_48 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_48;

architecture SYN_Behavioral of or2_48 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_47 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_47;

architecture SYN_Behavioral of or2_47 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_46 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_46;

architecture SYN_Behavioral of or2_46 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_45 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_45;

architecture SYN_Behavioral of or2_45 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_44 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_44;

architecture SYN_Behavioral of or2_44 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_43 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_43;

architecture SYN_Behavioral of or2_43 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_42 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_42;

architecture SYN_Behavioral of or2_42 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_41 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_41;

architecture SYN_Behavioral of or2_41 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_40 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_40;

architecture SYN_Behavioral of or2_40 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_39 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_39;

architecture SYN_Behavioral of or2_39 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_38 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_38;

architecture SYN_Behavioral of or2_38 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_37 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_37;

architecture SYN_Behavioral of or2_37 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_36 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_36;

architecture SYN_Behavioral of or2_36 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_35 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_35;

architecture SYN_Behavioral of or2_35 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_34 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_34;

architecture SYN_Behavioral of or2_34 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_33 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_33;

architecture SYN_Behavioral of or2_33 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_32 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_32;

architecture SYN_Behavioral of or2_32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_31 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_31;

architecture SYN_Behavioral of or2_31 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_30 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_30;

architecture SYN_Behavioral of or2_30 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_29 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_29;

architecture SYN_Behavioral of or2_29 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_28 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_28;

architecture SYN_Behavioral of or2_28 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_27 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_27;

architecture SYN_Behavioral of or2_27 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_26 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_26;

architecture SYN_Behavioral of or2_26 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_25 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_25;

architecture SYN_Behavioral of or2_25 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_24 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_24;

architecture SYN_Behavioral of or2_24 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_23 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_23;

architecture SYN_Behavioral of or2_23 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_22 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_22;

architecture SYN_Behavioral of or2_22 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_21 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_21;

architecture SYN_Behavioral of or2_21 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_20 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_20;

architecture SYN_Behavioral of or2_20 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_19 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_19;

architecture SYN_Behavioral of or2_19 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_18 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_18;

architecture SYN_Behavioral of or2_18 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_17 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_17;

architecture SYN_Behavioral of or2_17 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_16 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_16;

architecture SYN_Behavioral of or2_16 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_15 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_15;

architecture SYN_Behavioral of or2_15 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_14 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_14;

architecture SYN_Behavioral of or2_14 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_13 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_13;

architecture SYN_Behavioral of or2_13 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_12 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_12;

architecture SYN_Behavioral of or2_12 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_11 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_11;

architecture SYN_Behavioral of or2_11 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_10 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_10;

architecture SYN_Behavioral of or2_10 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_9 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_9;

architecture SYN_Behavioral of or2_9 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_8 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_8;

architecture SYN_Behavioral of or2_8 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_7 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_7;

architecture SYN_Behavioral of or2_7 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_6 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_6;

architecture SYN_Behavioral of or2_6 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_5 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_5;

architecture SYN_Behavioral of or2_5 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_4 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_4;

architecture SYN_Behavioral of or2_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_3 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_3;

architecture SYN_Behavioral of or2_3 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_2 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_2;

architecture SYN_Behavioral of or2_2 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_1 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_1;

architecture SYN_Behavioral of or2_1 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_440 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_440;

architecture SYN_Behavioral of xor2_440 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_439 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_439;

architecture SYN_Behavioral of xor2_439 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_438 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_438;

architecture SYN_Behavioral of xor2_438 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_437 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_437;

architecture SYN_Behavioral of xor2_437 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_436 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_436;

architecture SYN_Behavioral of xor2_436 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_435 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_435;

architecture SYN_Behavioral of xor2_435 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_434 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_434;

architecture SYN_Behavioral of xor2_434 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_433 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_433;

architecture SYN_Behavioral of xor2_433 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_432 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_432;

architecture SYN_Behavioral of xor2_432 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_431 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_431;

architecture SYN_Behavioral of xor2_431 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_430 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_430;

architecture SYN_Behavioral of xor2_430 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_429 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_429;

architecture SYN_Behavioral of xor2_429 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_428 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_428;

architecture SYN_Behavioral of xor2_428 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_427 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_427;

architecture SYN_Behavioral of xor2_427 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_426 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_426;

architecture SYN_Behavioral of xor2_426 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_425 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_425;

architecture SYN_Behavioral of xor2_425 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_424 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_424;

architecture SYN_Behavioral of xor2_424 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_423 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_423;

architecture SYN_Behavioral of xor2_423 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_422 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_422;

architecture SYN_Behavioral of xor2_422 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_421 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_421;

architecture SYN_Behavioral of xor2_421 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_420 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_420;

architecture SYN_Behavioral of xor2_420 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_419 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_419;

architecture SYN_Behavioral of xor2_419 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_418 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_418;

architecture SYN_Behavioral of xor2_418 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_417 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_417;

architecture SYN_Behavioral of xor2_417 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_416 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_416;

architecture SYN_Behavioral of xor2_416 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_415 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_415;

architecture SYN_Behavioral of xor2_415 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_414 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_414;

architecture SYN_Behavioral of xor2_414 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_413 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_413;

architecture SYN_Behavioral of xor2_413 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_412 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_412;

architecture SYN_Behavioral of xor2_412 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_411 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_411;

architecture SYN_Behavioral of xor2_411 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_410 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_410;

architecture SYN_Behavioral of xor2_410 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_409 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_409;

architecture SYN_Behavioral of xor2_409 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_408 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_408;

architecture SYN_Behavioral of xor2_408 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_407 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_407;

architecture SYN_Behavioral of xor2_407 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_406 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_406;

architecture SYN_Behavioral of xor2_406 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_405 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_405;

architecture SYN_Behavioral of xor2_405 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_404 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_404;

architecture SYN_Behavioral of xor2_404 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_403 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_403;

architecture SYN_Behavioral of xor2_403 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_402 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_402;

architecture SYN_Behavioral of xor2_402 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_401 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_401;

architecture SYN_Behavioral of xor2_401 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_400 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_400;

architecture SYN_Behavioral of xor2_400 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_399 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_399;

architecture SYN_Behavioral of xor2_399 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_398 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_398;

architecture SYN_Behavioral of xor2_398 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_397 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_397;

architecture SYN_Behavioral of xor2_397 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_396 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_396;

architecture SYN_Behavioral of xor2_396 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_395 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_395;

architecture SYN_Behavioral of xor2_395 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_394 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_394;

architecture SYN_Behavioral of xor2_394 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_393 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_393;

architecture SYN_Behavioral of xor2_393 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_392 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_392;

architecture SYN_Behavioral of xor2_392 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_391 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_391;

architecture SYN_Behavioral of xor2_391 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_390 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_390;

architecture SYN_Behavioral of xor2_390 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_389 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_389;

architecture SYN_Behavioral of xor2_389 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_388 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_388;

architecture SYN_Behavioral of xor2_388 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_387 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_387;

architecture SYN_Behavioral of xor2_387 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_386 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_386;

architecture SYN_Behavioral of xor2_386 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_385 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_385;

architecture SYN_Behavioral of xor2_385 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_384 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_384;

architecture SYN_Behavioral of xor2_384 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_383 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_383;

architecture SYN_Behavioral of xor2_383 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_382 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_382;

architecture SYN_Behavioral of xor2_382 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_381 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_381;

architecture SYN_Behavioral of xor2_381 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_380 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_380;

architecture SYN_Behavioral of xor2_380 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_379 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_379;

architecture SYN_Behavioral of xor2_379 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_378 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_378;

architecture SYN_Behavioral of xor2_378 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_377 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_377;

architecture SYN_Behavioral of xor2_377 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_376 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_376;

architecture SYN_Behavioral of xor2_376 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_375 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_375;

architecture SYN_Behavioral of xor2_375 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_374 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_374;

architecture SYN_Behavioral of xor2_374 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_373 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_373;

architecture SYN_Behavioral of xor2_373 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_372 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_372;

architecture SYN_Behavioral of xor2_372 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_371 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_371;

architecture SYN_Behavioral of xor2_371 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_370 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_370;

architecture SYN_Behavioral of xor2_370 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_369 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_369;

architecture SYN_Behavioral of xor2_369 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_368 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_368;

architecture SYN_Behavioral of xor2_368 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_367 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_367;

architecture SYN_Behavioral of xor2_367 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_366 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_366;

architecture SYN_Behavioral of xor2_366 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_365 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_365;

architecture SYN_Behavioral of xor2_365 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_364 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_364;

architecture SYN_Behavioral of xor2_364 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_363 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_363;

architecture SYN_Behavioral of xor2_363 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_362 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_362;

architecture SYN_Behavioral of xor2_362 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_361 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_361;

architecture SYN_Behavioral of xor2_361 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_360 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_360;

architecture SYN_Behavioral of xor2_360 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_359 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_359;

architecture SYN_Behavioral of xor2_359 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_358 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_358;

architecture SYN_Behavioral of xor2_358 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_357 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_357;

architecture SYN_Behavioral of xor2_357 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_356 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_356;

architecture SYN_Behavioral of xor2_356 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_355 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_355;

architecture SYN_Behavioral of xor2_355 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_354 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_354;

architecture SYN_Behavioral of xor2_354 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_353 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_353;

architecture SYN_Behavioral of xor2_353 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_352 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_352;

architecture SYN_Behavioral of xor2_352 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_351 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_351;

architecture SYN_Behavioral of xor2_351 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_350 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_350;

architecture SYN_Behavioral of xor2_350 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_349 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_349;

architecture SYN_Behavioral of xor2_349 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_348 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_348;

architecture SYN_Behavioral of xor2_348 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_347 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_347;

architecture SYN_Behavioral of xor2_347 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_346 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_346;

architecture SYN_Behavioral of xor2_346 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_345 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_345;

architecture SYN_Behavioral of xor2_345 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_344 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_344;

architecture SYN_Behavioral of xor2_344 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_343 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_343;

architecture SYN_Behavioral of xor2_343 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_342 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_342;

architecture SYN_Behavioral of xor2_342 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_341 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_341;

architecture SYN_Behavioral of xor2_341 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_340 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_340;

architecture SYN_Behavioral of xor2_340 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_339 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_339;

architecture SYN_Behavioral of xor2_339 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_338 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_338;

architecture SYN_Behavioral of xor2_338 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_337 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_337;

architecture SYN_Behavioral of xor2_337 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_336 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_336;

architecture SYN_Behavioral of xor2_336 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_335 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_335;

architecture SYN_Behavioral of xor2_335 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_334 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_334;

architecture SYN_Behavioral of xor2_334 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_333 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_333;

architecture SYN_Behavioral of xor2_333 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_332 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_332;

architecture SYN_Behavioral of xor2_332 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_331 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_331;

architecture SYN_Behavioral of xor2_331 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_330 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_330;

architecture SYN_Behavioral of xor2_330 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_329 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_329;

architecture SYN_Behavioral of xor2_329 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_328 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_328;

architecture SYN_Behavioral of xor2_328 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_327 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_327;

architecture SYN_Behavioral of xor2_327 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_326 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_326;

architecture SYN_Behavioral of xor2_326 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_325 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_325;

architecture SYN_Behavioral of xor2_325 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_324 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_324;

architecture SYN_Behavioral of xor2_324 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_323 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_323;

architecture SYN_Behavioral of xor2_323 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_322 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_322;

architecture SYN_Behavioral of xor2_322 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_321 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_321;

architecture SYN_Behavioral of xor2_321 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_320 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_320;

architecture SYN_Behavioral of xor2_320 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_319 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_319;

architecture SYN_Behavioral of xor2_319 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_318 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_318;

architecture SYN_Behavioral of xor2_318 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_317 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_317;

architecture SYN_Behavioral of xor2_317 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_316 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_316;

architecture SYN_Behavioral of xor2_316 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_315 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_315;

architecture SYN_Behavioral of xor2_315 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_314 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_314;

architecture SYN_Behavioral of xor2_314 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_313 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_313;

architecture SYN_Behavioral of xor2_313 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_312 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_312;

architecture SYN_Behavioral of xor2_312 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_311 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_311;

architecture SYN_Behavioral of xor2_311 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_310 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_310;

architecture SYN_Behavioral of xor2_310 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_309 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_309;

architecture SYN_Behavioral of xor2_309 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_308 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_308;

architecture SYN_Behavioral of xor2_308 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_307 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_307;

architecture SYN_Behavioral of xor2_307 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_306 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_306;

architecture SYN_Behavioral of xor2_306 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_305 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_305;

architecture SYN_Behavioral of xor2_305 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_304 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_304;

architecture SYN_Behavioral of xor2_304 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_303 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_303;

architecture SYN_Behavioral of xor2_303 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_302 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_302;

architecture SYN_Behavioral of xor2_302 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_301 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_301;

architecture SYN_Behavioral of xor2_301 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_300 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_300;

architecture SYN_Behavioral of xor2_300 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_299 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_299;

architecture SYN_Behavioral of xor2_299 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_298 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_298;

architecture SYN_Behavioral of xor2_298 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_297 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_297;

architecture SYN_Behavioral of xor2_297 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_296 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_296;

architecture SYN_Behavioral of xor2_296 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_295 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_295;

architecture SYN_Behavioral of xor2_295 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_294 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_294;

architecture SYN_Behavioral of xor2_294 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_293 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_293;

architecture SYN_Behavioral of xor2_293 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_292 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_292;

architecture SYN_Behavioral of xor2_292 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_291 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_291;

architecture SYN_Behavioral of xor2_291 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_290 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_290;

architecture SYN_Behavioral of xor2_290 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_289 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_289;

architecture SYN_Behavioral of xor2_289 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_288 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_288;

architecture SYN_Behavioral of xor2_288 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_287 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_287;

architecture SYN_Behavioral of xor2_287 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_286 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_286;

architecture SYN_Behavioral of xor2_286 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_285 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_285;

architecture SYN_Behavioral of xor2_285 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_284 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_284;

architecture SYN_Behavioral of xor2_284 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_283 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_283;

architecture SYN_Behavioral of xor2_283 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_282 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_282;

architecture SYN_Behavioral of xor2_282 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_281 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_281;

architecture SYN_Behavioral of xor2_281 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_280 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_280;

architecture SYN_Behavioral of xor2_280 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_279 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_279;

architecture SYN_Behavioral of xor2_279 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_278 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_278;

architecture SYN_Behavioral of xor2_278 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_277 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_277;

architecture SYN_Behavioral of xor2_277 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_276 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_276;

architecture SYN_Behavioral of xor2_276 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_275 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_275;

architecture SYN_Behavioral of xor2_275 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_274 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_274;

architecture SYN_Behavioral of xor2_274 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_273 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_273;

architecture SYN_Behavioral of xor2_273 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_272 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_272;

architecture SYN_Behavioral of xor2_272 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_271 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_271;

architecture SYN_Behavioral of xor2_271 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_270 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_270;

architecture SYN_Behavioral of xor2_270 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_269 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_269;

architecture SYN_Behavioral of xor2_269 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_268 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_268;

architecture SYN_Behavioral of xor2_268 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_267 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_267;

architecture SYN_Behavioral of xor2_267 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_266 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_266;

architecture SYN_Behavioral of xor2_266 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_265 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_265;

architecture SYN_Behavioral of xor2_265 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_264 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_264;

architecture SYN_Behavioral of xor2_264 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_263 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_263;

architecture SYN_Behavioral of xor2_263 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_262 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_262;

architecture SYN_Behavioral of xor2_262 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_261 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_261;

architecture SYN_Behavioral of xor2_261 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_260 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_260;

architecture SYN_Behavioral of xor2_260 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_259 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_259;

architecture SYN_Behavioral of xor2_259 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_258 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_258;

architecture SYN_Behavioral of xor2_258 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_257 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_257;

architecture SYN_Behavioral of xor2_257 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_256 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_256;

architecture SYN_Behavioral of xor2_256 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_255 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_255;

architecture SYN_Behavioral of xor2_255 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_254 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_254;

architecture SYN_Behavioral of xor2_254 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_253 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_253;

architecture SYN_Behavioral of xor2_253 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_252 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_252;

architecture SYN_Behavioral of xor2_252 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_251 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_251;

architecture SYN_Behavioral of xor2_251 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_250 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_250;

architecture SYN_Behavioral of xor2_250 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_249 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_249;

architecture SYN_Behavioral of xor2_249 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_248 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_248;

architecture SYN_Behavioral of xor2_248 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_247 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_247;

architecture SYN_Behavioral of xor2_247 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_246 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_246;

architecture SYN_Behavioral of xor2_246 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_245 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_245;

architecture SYN_Behavioral of xor2_245 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_244 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_244;

architecture SYN_Behavioral of xor2_244 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_243 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_243;

architecture SYN_Behavioral of xor2_243 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_242 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_242;

architecture SYN_Behavioral of xor2_242 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_241 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_241;

architecture SYN_Behavioral of xor2_241 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_240 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_240;

architecture SYN_Behavioral of xor2_240 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_239 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_239;

architecture SYN_Behavioral of xor2_239 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_238 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_238;

architecture SYN_Behavioral of xor2_238 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_237 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_237;

architecture SYN_Behavioral of xor2_237 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_236 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_236;

architecture SYN_Behavioral of xor2_236 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_235 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_235;

architecture SYN_Behavioral of xor2_235 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_234 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_234;

architecture SYN_Behavioral of xor2_234 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_233 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_233;

architecture SYN_Behavioral of xor2_233 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_232 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_232;

architecture SYN_Behavioral of xor2_232 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_231 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_231;

architecture SYN_Behavioral of xor2_231 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_230 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_230;

architecture SYN_Behavioral of xor2_230 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_229 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_229;

architecture SYN_Behavioral of xor2_229 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_228 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_228;

architecture SYN_Behavioral of xor2_228 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_227 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_227;

architecture SYN_Behavioral of xor2_227 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_226 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_226;

architecture SYN_Behavioral of xor2_226 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_225 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_225;

architecture SYN_Behavioral of xor2_225 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_224 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_224;

architecture SYN_Behavioral of xor2_224 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_223 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_223;

architecture SYN_Behavioral of xor2_223 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_222 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_222;

architecture SYN_Behavioral of xor2_222 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_221 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_221;

architecture SYN_Behavioral of xor2_221 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_220 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_220;

architecture SYN_Behavioral of xor2_220 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_219 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_219;

architecture SYN_Behavioral of xor2_219 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_218 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_218;

architecture SYN_Behavioral of xor2_218 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_217 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_217;

architecture SYN_Behavioral of xor2_217 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_216 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_216;

architecture SYN_Behavioral of xor2_216 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_215 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_215;

architecture SYN_Behavioral of xor2_215 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_214 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_214;

architecture SYN_Behavioral of xor2_214 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_213 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_213;

architecture SYN_Behavioral of xor2_213 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_212 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_212;

architecture SYN_Behavioral of xor2_212 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_211 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_211;

architecture SYN_Behavioral of xor2_211 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_210 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_210;

architecture SYN_Behavioral of xor2_210 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_209 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_209;

architecture SYN_Behavioral of xor2_209 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_208 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_208;

architecture SYN_Behavioral of xor2_208 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_207 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_207;

architecture SYN_Behavioral of xor2_207 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_206 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_206;

architecture SYN_Behavioral of xor2_206 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_205 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_205;

architecture SYN_Behavioral of xor2_205 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_204 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_204;

architecture SYN_Behavioral of xor2_204 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_203 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_203;

architecture SYN_Behavioral of xor2_203 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_202 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_202;

architecture SYN_Behavioral of xor2_202 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_201 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_201;

architecture SYN_Behavioral of xor2_201 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_200 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_200;

architecture SYN_Behavioral of xor2_200 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_199 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_199;

architecture SYN_Behavioral of xor2_199 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_198 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_198;

architecture SYN_Behavioral of xor2_198 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_197 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_197;

architecture SYN_Behavioral of xor2_197 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_196 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_196;

architecture SYN_Behavioral of xor2_196 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_195 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_195;

architecture SYN_Behavioral of xor2_195 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_194 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_194;

architecture SYN_Behavioral of xor2_194 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_193 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_193;

architecture SYN_Behavioral of xor2_193 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_192 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_192;

architecture SYN_Behavioral of xor2_192 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_191 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_191;

architecture SYN_Behavioral of xor2_191 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_190 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_190;

architecture SYN_Behavioral of xor2_190 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_189 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_189;

architecture SYN_Behavioral of xor2_189 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_188 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_188;

architecture SYN_Behavioral of xor2_188 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_187 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_187;

architecture SYN_Behavioral of xor2_187 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_186 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_186;

architecture SYN_Behavioral of xor2_186 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_185 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_185;

architecture SYN_Behavioral of xor2_185 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_184 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_184;

architecture SYN_Behavioral of xor2_184 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_183 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_183;

architecture SYN_Behavioral of xor2_183 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_182 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_182;

architecture SYN_Behavioral of xor2_182 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_181 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_181;

architecture SYN_Behavioral of xor2_181 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_180 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_180;

architecture SYN_Behavioral of xor2_180 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_179 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_179;

architecture SYN_Behavioral of xor2_179 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_178 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_178;

architecture SYN_Behavioral of xor2_178 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_177 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_177;

architecture SYN_Behavioral of xor2_177 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_176 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_176;

architecture SYN_Behavioral of xor2_176 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_175 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_175;

architecture SYN_Behavioral of xor2_175 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_174 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_174;

architecture SYN_Behavioral of xor2_174 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_173 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_173;

architecture SYN_Behavioral of xor2_173 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_172 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_172;

architecture SYN_Behavioral of xor2_172 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_171 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_171;

architecture SYN_Behavioral of xor2_171 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_170 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_170;

architecture SYN_Behavioral of xor2_170 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_169 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_169;

architecture SYN_Behavioral of xor2_169 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_168 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_168;

architecture SYN_Behavioral of xor2_168 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_167 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_167;

architecture SYN_Behavioral of xor2_167 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_166 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_166;

architecture SYN_Behavioral of xor2_166 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_165 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_165;

architecture SYN_Behavioral of xor2_165 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_164 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_164;

architecture SYN_Behavioral of xor2_164 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_163 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_163;

architecture SYN_Behavioral of xor2_163 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_162 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_162;

architecture SYN_Behavioral of xor2_162 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_161 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_161;

architecture SYN_Behavioral of xor2_161 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_160 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_160;

architecture SYN_Behavioral of xor2_160 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_159 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_159;

architecture SYN_Behavioral of xor2_159 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_158 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_158;

architecture SYN_Behavioral of xor2_158 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_157 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_157;

architecture SYN_Behavioral of xor2_157 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_156 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_156;

architecture SYN_Behavioral of xor2_156 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_155 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_155;

architecture SYN_Behavioral of xor2_155 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_154 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_154;

architecture SYN_Behavioral of xor2_154 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_153 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_153;

architecture SYN_Behavioral of xor2_153 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_152 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_152;

architecture SYN_Behavioral of xor2_152 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_151 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_151;

architecture SYN_Behavioral of xor2_151 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_150 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_150;

architecture SYN_Behavioral of xor2_150 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_149 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_149;

architecture SYN_Behavioral of xor2_149 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_148 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_148;

architecture SYN_Behavioral of xor2_148 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_147 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_147;

architecture SYN_Behavioral of xor2_147 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_146 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_146;

architecture SYN_Behavioral of xor2_146 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_145 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_145;

architecture SYN_Behavioral of xor2_145 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_144 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_144;

architecture SYN_Behavioral of xor2_144 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_143 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_143;

architecture SYN_Behavioral of xor2_143 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_142 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_142;

architecture SYN_Behavioral of xor2_142 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_141 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_141;

architecture SYN_Behavioral of xor2_141 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_140 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_140;

architecture SYN_Behavioral of xor2_140 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_139 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_139;

architecture SYN_Behavioral of xor2_139 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_138 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_138;

architecture SYN_Behavioral of xor2_138 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_137 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_137;

architecture SYN_Behavioral of xor2_137 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_136 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_136;

architecture SYN_Behavioral of xor2_136 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_135 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_135;

architecture SYN_Behavioral of xor2_135 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_134 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_134;

architecture SYN_Behavioral of xor2_134 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_133 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_133;

architecture SYN_Behavioral of xor2_133 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_132 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_132;

architecture SYN_Behavioral of xor2_132 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_131 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_131;

architecture SYN_Behavioral of xor2_131 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_130 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_130;

architecture SYN_Behavioral of xor2_130 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_129 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_129;

architecture SYN_Behavioral of xor2_129 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_128 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_128;

architecture SYN_Behavioral of xor2_128 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_127 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_127;

architecture SYN_Behavioral of xor2_127 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_126 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_126;

architecture SYN_Behavioral of xor2_126 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_125 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_125;

architecture SYN_Behavioral of xor2_125 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_124 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_124;

architecture SYN_Behavioral of xor2_124 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_123 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_123;

architecture SYN_Behavioral of xor2_123 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_122 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_122;

architecture SYN_Behavioral of xor2_122 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_121 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_121;

architecture SYN_Behavioral of xor2_121 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_120 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_120;

architecture SYN_Behavioral of xor2_120 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_119 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_119;

architecture SYN_Behavioral of xor2_119 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_118 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_118;

architecture SYN_Behavioral of xor2_118 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_117 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_117;

architecture SYN_Behavioral of xor2_117 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_116 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_116;

architecture SYN_Behavioral of xor2_116 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_115 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_115;

architecture SYN_Behavioral of xor2_115 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_114 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_114;

architecture SYN_Behavioral of xor2_114 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_113 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_113;

architecture SYN_Behavioral of xor2_113 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_112 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_112;

architecture SYN_Behavioral of xor2_112 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_111 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_111;

architecture SYN_Behavioral of xor2_111 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_110 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_110;

architecture SYN_Behavioral of xor2_110 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_109 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_109;

architecture SYN_Behavioral of xor2_109 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_108 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_108;

architecture SYN_Behavioral of xor2_108 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_107 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_107;

architecture SYN_Behavioral of xor2_107 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_106 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_106;

architecture SYN_Behavioral of xor2_106 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_105 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_105;

architecture SYN_Behavioral of xor2_105 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_104 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_104;

architecture SYN_Behavioral of xor2_104 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_103 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_103;

architecture SYN_Behavioral of xor2_103 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_102 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_102;

architecture SYN_Behavioral of xor2_102 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_101 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_101;

architecture SYN_Behavioral of xor2_101 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_100 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_100;

architecture SYN_Behavioral of xor2_100 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_99 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_99;

architecture SYN_Behavioral of xor2_99 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_98 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_98;

architecture SYN_Behavioral of xor2_98 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_97 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_97;

architecture SYN_Behavioral of xor2_97 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_96 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_96;

architecture SYN_Behavioral of xor2_96 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_95 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_95;

architecture SYN_Behavioral of xor2_95 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_94 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_94;

architecture SYN_Behavioral of xor2_94 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_93 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_93;

architecture SYN_Behavioral of xor2_93 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_92 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_92;

architecture SYN_Behavioral of xor2_92 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_91 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_91;

architecture SYN_Behavioral of xor2_91 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_90 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_90;

architecture SYN_Behavioral of xor2_90 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_89 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_89;

architecture SYN_Behavioral of xor2_89 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_88 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_88;

architecture SYN_Behavioral of xor2_88 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_87 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_87;

architecture SYN_Behavioral of xor2_87 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_86 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_86;

architecture SYN_Behavioral of xor2_86 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_85 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_85;

architecture SYN_Behavioral of xor2_85 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_84 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_84;

architecture SYN_Behavioral of xor2_84 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_83 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_83;

architecture SYN_Behavioral of xor2_83 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_82 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_82;

architecture SYN_Behavioral of xor2_82 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_81 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_81;

architecture SYN_Behavioral of xor2_81 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_80 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_80;

architecture SYN_Behavioral of xor2_80 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_79 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_79;

architecture SYN_Behavioral of xor2_79 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_78 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_78;

architecture SYN_Behavioral of xor2_78 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_77 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_77;

architecture SYN_Behavioral of xor2_77 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_76 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_76;

architecture SYN_Behavioral of xor2_76 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_75 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_75;

architecture SYN_Behavioral of xor2_75 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_74 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_74;

architecture SYN_Behavioral of xor2_74 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_73 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_73;

architecture SYN_Behavioral of xor2_73 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_72 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_72;

architecture SYN_Behavioral of xor2_72 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_71 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_71;

architecture SYN_Behavioral of xor2_71 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_70 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_70;

architecture SYN_Behavioral of xor2_70 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_69 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_69;

architecture SYN_Behavioral of xor2_69 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_68 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_68;

architecture SYN_Behavioral of xor2_68 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_67 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_67;

architecture SYN_Behavioral of xor2_67 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_66 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_66;

architecture SYN_Behavioral of xor2_66 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_65 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_65;

architecture SYN_Behavioral of xor2_65 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_64 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_64;

architecture SYN_Behavioral of xor2_64 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_63 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_63;

architecture SYN_Behavioral of xor2_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_62 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_62;

architecture SYN_Behavioral of xor2_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_61 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_61;

architecture SYN_Behavioral of xor2_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_60 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_60;

architecture SYN_Behavioral of xor2_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_59 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_59;

architecture SYN_Behavioral of xor2_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_58 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_58;

architecture SYN_Behavioral of xor2_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_57 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_57;

architecture SYN_Behavioral of xor2_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_56 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_56;

architecture SYN_Behavioral of xor2_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_55 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_55;

architecture SYN_Behavioral of xor2_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_54 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_54;

architecture SYN_Behavioral of xor2_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_53 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_53;

architecture SYN_Behavioral of xor2_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_52 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_52;

architecture SYN_Behavioral of xor2_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_51 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_51;

architecture SYN_Behavioral of xor2_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_50 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_50;

architecture SYN_Behavioral of xor2_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_49 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_49;

architecture SYN_Behavioral of xor2_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_48 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_48;

architecture SYN_Behavioral of xor2_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_47 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_47;

architecture SYN_Behavioral of xor2_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_46 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_46;

architecture SYN_Behavioral of xor2_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_45 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_45;

architecture SYN_Behavioral of xor2_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_44 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_44;

architecture SYN_Behavioral of xor2_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_43 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_43;

architecture SYN_Behavioral of xor2_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_42 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_42;

architecture SYN_Behavioral of xor2_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_41 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_41;

architecture SYN_Behavioral of xor2_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_40 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_40;

architecture SYN_Behavioral of xor2_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_39 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_39;

architecture SYN_Behavioral of xor2_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_38 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_38;

architecture SYN_Behavioral of xor2_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_37 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_37;

architecture SYN_Behavioral of xor2_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_36 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_36;

architecture SYN_Behavioral of xor2_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_35 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_35;

architecture SYN_Behavioral of xor2_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_34 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_34;

architecture SYN_Behavioral of xor2_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_33 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_33;

architecture SYN_Behavioral of xor2_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_32 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_32;

architecture SYN_Behavioral of xor2_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_31 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_31;

architecture SYN_Behavioral of xor2_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_30 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_30;

architecture SYN_Behavioral of xor2_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_29 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_29;

architecture SYN_Behavioral of xor2_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_28 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_28;

architecture SYN_Behavioral of xor2_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_27 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_27;

architecture SYN_Behavioral of xor2_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_26 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_26;

architecture SYN_Behavioral of xor2_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_25 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_25;

architecture SYN_Behavioral of xor2_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_24 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_24;

architecture SYN_Behavioral of xor2_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_23 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_23;

architecture SYN_Behavioral of xor2_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_22 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_22;

architecture SYN_Behavioral of xor2_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_21 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_21;

architecture SYN_Behavioral of xor2_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_20 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_20;

architecture SYN_Behavioral of xor2_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_19 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_19;

architecture SYN_Behavioral of xor2_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_18 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_18;

architecture SYN_Behavioral of xor2_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_17 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_17;

architecture SYN_Behavioral of xor2_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_16 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_16;

architecture SYN_Behavioral of xor2_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_15 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_15;

architecture SYN_Behavioral of xor2_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_14 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_14;

architecture SYN_Behavioral of xor2_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_13 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_13;

architecture SYN_Behavioral of xor2_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_12 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_12;

architecture SYN_Behavioral of xor2_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_11 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_11;

architecture SYN_Behavioral of xor2_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_10 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_10;

architecture SYN_Behavioral of xor2_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_9 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_9;

architecture SYN_Behavioral of xor2_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_8 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_8;

architecture SYN_Behavioral of xor2_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_7 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_7;

architecture SYN_Behavioral of xor2_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_6 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_6;

architecture SYN_Behavioral of xor2_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_5 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_5;

architecture SYN_Behavioral of xor2_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_4 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_4;

architecture SYN_Behavioral of xor2_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_3 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_3;

architecture SYN_Behavioral of xor2_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_2 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_2;

architecture SYN_Behavioral of xor2_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_1 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_1;

architecture SYN_Behavioral of xor2_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_440 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_440;

architecture SYN_Behavioral of and2_440 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_439 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_439;

architecture SYN_Behavioral of and2_439 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_438 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_438;

architecture SYN_Behavioral of and2_438 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_437 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_437;

architecture SYN_Behavioral of and2_437 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_436 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_436;

architecture SYN_Behavioral of and2_436 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_435 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_435;

architecture SYN_Behavioral of and2_435 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_434 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_434;

architecture SYN_Behavioral of and2_434 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_433 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_433;

architecture SYN_Behavioral of and2_433 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_432 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_432;

architecture SYN_Behavioral of and2_432 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_431 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_431;

architecture SYN_Behavioral of and2_431 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_430 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_430;

architecture SYN_Behavioral of and2_430 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_429 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_429;

architecture SYN_Behavioral of and2_429 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_428 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_428;

architecture SYN_Behavioral of and2_428 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_427 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_427;

architecture SYN_Behavioral of and2_427 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_426 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_426;

architecture SYN_Behavioral of and2_426 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_425 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_425;

architecture SYN_Behavioral of and2_425 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_424 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_424;

architecture SYN_Behavioral of and2_424 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_423 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_423;

architecture SYN_Behavioral of and2_423 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_422 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_422;

architecture SYN_Behavioral of and2_422 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_421 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_421;

architecture SYN_Behavioral of and2_421 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_420 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_420;

architecture SYN_Behavioral of and2_420 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_419 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_419;

architecture SYN_Behavioral of and2_419 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_418 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_418;

architecture SYN_Behavioral of and2_418 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_417 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_417;

architecture SYN_Behavioral of and2_417 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_416 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_416;

architecture SYN_Behavioral of and2_416 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_415 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_415;

architecture SYN_Behavioral of and2_415 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_414 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_414;

architecture SYN_Behavioral of and2_414 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_413 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_413;

architecture SYN_Behavioral of and2_413 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_412 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_412;

architecture SYN_Behavioral of and2_412 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_411 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_411;

architecture SYN_Behavioral of and2_411 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_410 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_410;

architecture SYN_Behavioral of and2_410 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_409 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_409;

architecture SYN_Behavioral of and2_409 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_408 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_408;

architecture SYN_Behavioral of and2_408 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_407 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_407;

architecture SYN_Behavioral of and2_407 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_406 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_406;

architecture SYN_Behavioral of and2_406 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_405 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_405;

architecture SYN_Behavioral of and2_405 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_404 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_404;

architecture SYN_Behavioral of and2_404 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_403 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_403;

architecture SYN_Behavioral of and2_403 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_402 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_402;

architecture SYN_Behavioral of and2_402 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_401 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_401;

architecture SYN_Behavioral of and2_401 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_400 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_400;

architecture SYN_Behavioral of and2_400 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_399 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_399;

architecture SYN_Behavioral of and2_399 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_398 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_398;

architecture SYN_Behavioral of and2_398 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_397 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_397;

architecture SYN_Behavioral of and2_397 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_396 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_396;

architecture SYN_Behavioral of and2_396 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_395 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_395;

architecture SYN_Behavioral of and2_395 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_394 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_394;

architecture SYN_Behavioral of and2_394 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_393 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_393;

architecture SYN_Behavioral of and2_393 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_392 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_392;

architecture SYN_Behavioral of and2_392 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_391 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_391;

architecture SYN_Behavioral of and2_391 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_390 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_390;

architecture SYN_Behavioral of and2_390 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_389 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_389;

architecture SYN_Behavioral of and2_389 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_388 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_388;

architecture SYN_Behavioral of and2_388 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_387 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_387;

architecture SYN_Behavioral of and2_387 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_386 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_386;

architecture SYN_Behavioral of and2_386 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_385 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_385;

architecture SYN_Behavioral of and2_385 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_384 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_384;

architecture SYN_Behavioral of and2_384 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_383 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_383;

architecture SYN_Behavioral of and2_383 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_382 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_382;

architecture SYN_Behavioral of and2_382 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_381 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_381;

architecture SYN_Behavioral of and2_381 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_380 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_380;

architecture SYN_Behavioral of and2_380 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_379 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_379;

architecture SYN_Behavioral of and2_379 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_378 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_378;

architecture SYN_Behavioral of and2_378 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_377 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_377;

architecture SYN_Behavioral of and2_377 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_376 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_376;

architecture SYN_Behavioral of and2_376 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_375 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_375;

architecture SYN_Behavioral of and2_375 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_374 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_374;

architecture SYN_Behavioral of and2_374 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_373 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_373;

architecture SYN_Behavioral of and2_373 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_372 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_372;

architecture SYN_Behavioral of and2_372 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_371 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_371;

architecture SYN_Behavioral of and2_371 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_370 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_370;

architecture SYN_Behavioral of and2_370 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_369 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_369;

architecture SYN_Behavioral of and2_369 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_368 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_368;

architecture SYN_Behavioral of and2_368 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_367 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_367;

architecture SYN_Behavioral of and2_367 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_366 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_366;

architecture SYN_Behavioral of and2_366 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_365 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_365;

architecture SYN_Behavioral of and2_365 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_364 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_364;

architecture SYN_Behavioral of and2_364 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_363 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_363;

architecture SYN_Behavioral of and2_363 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_362 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_362;

architecture SYN_Behavioral of and2_362 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_361 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_361;

architecture SYN_Behavioral of and2_361 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_360 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_360;

architecture SYN_Behavioral of and2_360 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_359 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_359;

architecture SYN_Behavioral of and2_359 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_358 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_358;

architecture SYN_Behavioral of and2_358 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_357 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_357;

architecture SYN_Behavioral of and2_357 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_356 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_356;

architecture SYN_Behavioral of and2_356 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_355 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_355;

architecture SYN_Behavioral of and2_355 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_354 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_354;

architecture SYN_Behavioral of and2_354 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_353 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_353;

architecture SYN_Behavioral of and2_353 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_352 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_352;

architecture SYN_Behavioral of and2_352 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_351 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_351;

architecture SYN_Behavioral of and2_351 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_350 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_350;

architecture SYN_Behavioral of and2_350 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_349 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_349;

architecture SYN_Behavioral of and2_349 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_348 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_348;

architecture SYN_Behavioral of and2_348 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_347 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_347;

architecture SYN_Behavioral of and2_347 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_346 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_346;

architecture SYN_Behavioral of and2_346 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_345 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_345;

architecture SYN_Behavioral of and2_345 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_344 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_344;

architecture SYN_Behavioral of and2_344 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_343 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_343;

architecture SYN_Behavioral of and2_343 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_342 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_342;

architecture SYN_Behavioral of and2_342 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_341 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_341;

architecture SYN_Behavioral of and2_341 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_340 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_340;

architecture SYN_Behavioral of and2_340 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_339 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_339;

architecture SYN_Behavioral of and2_339 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_338 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_338;

architecture SYN_Behavioral of and2_338 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_337 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_337;

architecture SYN_Behavioral of and2_337 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_336 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_336;

architecture SYN_Behavioral of and2_336 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_335 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_335;

architecture SYN_Behavioral of and2_335 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_334 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_334;

architecture SYN_Behavioral of and2_334 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_333 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_333;

architecture SYN_Behavioral of and2_333 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_332 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_332;

architecture SYN_Behavioral of and2_332 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_331 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_331;

architecture SYN_Behavioral of and2_331 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_330 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_330;

architecture SYN_Behavioral of and2_330 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_329 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_329;

architecture SYN_Behavioral of and2_329 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_328 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_328;

architecture SYN_Behavioral of and2_328 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_327 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_327;

architecture SYN_Behavioral of and2_327 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_326 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_326;

architecture SYN_Behavioral of and2_326 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_325 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_325;

architecture SYN_Behavioral of and2_325 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_324 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_324;

architecture SYN_Behavioral of and2_324 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_323 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_323;

architecture SYN_Behavioral of and2_323 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_322 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_322;

architecture SYN_Behavioral of and2_322 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_321 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_321;

architecture SYN_Behavioral of and2_321 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_320 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_320;

architecture SYN_Behavioral of and2_320 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_319 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_319;

architecture SYN_Behavioral of and2_319 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_318 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_318;

architecture SYN_Behavioral of and2_318 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_317 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_317;

architecture SYN_Behavioral of and2_317 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_316 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_316;

architecture SYN_Behavioral of and2_316 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_315 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_315;

architecture SYN_Behavioral of and2_315 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_314 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_314;

architecture SYN_Behavioral of and2_314 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_313 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_313;

architecture SYN_Behavioral of and2_313 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_312 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_312;

architecture SYN_Behavioral of and2_312 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_311 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_311;

architecture SYN_Behavioral of and2_311 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_310 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_310;

architecture SYN_Behavioral of and2_310 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_309 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_309;

architecture SYN_Behavioral of and2_309 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_308 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_308;

architecture SYN_Behavioral of and2_308 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_307 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_307;

architecture SYN_Behavioral of and2_307 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_306 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_306;

architecture SYN_Behavioral of and2_306 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_305 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_305;

architecture SYN_Behavioral of and2_305 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_304 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_304;

architecture SYN_Behavioral of and2_304 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_303 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_303;

architecture SYN_Behavioral of and2_303 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_302 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_302;

architecture SYN_Behavioral of and2_302 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_301 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_301;

architecture SYN_Behavioral of and2_301 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_300 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_300;

architecture SYN_Behavioral of and2_300 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_299 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_299;

architecture SYN_Behavioral of and2_299 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_298 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_298;

architecture SYN_Behavioral of and2_298 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_297 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_297;

architecture SYN_Behavioral of and2_297 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_296 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_296;

architecture SYN_Behavioral of and2_296 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_295 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_295;

architecture SYN_Behavioral of and2_295 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_294 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_294;

architecture SYN_Behavioral of and2_294 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_293 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_293;

architecture SYN_Behavioral of and2_293 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_292 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_292;

architecture SYN_Behavioral of and2_292 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_291 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_291;

architecture SYN_Behavioral of and2_291 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_290 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_290;

architecture SYN_Behavioral of and2_290 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_289 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_289;

architecture SYN_Behavioral of and2_289 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_288 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_288;

architecture SYN_Behavioral of and2_288 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_287 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_287;

architecture SYN_Behavioral of and2_287 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_286 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_286;

architecture SYN_Behavioral of and2_286 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_285 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_285;

architecture SYN_Behavioral of and2_285 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_284 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_284;

architecture SYN_Behavioral of and2_284 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_283 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_283;

architecture SYN_Behavioral of and2_283 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_282 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_282;

architecture SYN_Behavioral of and2_282 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_281 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_281;

architecture SYN_Behavioral of and2_281 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_280 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_280;

architecture SYN_Behavioral of and2_280 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_279 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_279;

architecture SYN_Behavioral of and2_279 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_278 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_278;

architecture SYN_Behavioral of and2_278 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_277 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_277;

architecture SYN_Behavioral of and2_277 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_276 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_276;

architecture SYN_Behavioral of and2_276 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_275 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_275;

architecture SYN_Behavioral of and2_275 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_274 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_274;

architecture SYN_Behavioral of and2_274 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_273 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_273;

architecture SYN_Behavioral of and2_273 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_272 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_272;

architecture SYN_Behavioral of and2_272 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_271 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_271;

architecture SYN_Behavioral of and2_271 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_270 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_270;

architecture SYN_Behavioral of and2_270 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_269 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_269;

architecture SYN_Behavioral of and2_269 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_268 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_268;

architecture SYN_Behavioral of and2_268 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_267 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_267;

architecture SYN_Behavioral of and2_267 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_266 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_266;

architecture SYN_Behavioral of and2_266 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_265 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_265;

architecture SYN_Behavioral of and2_265 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_264 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_264;

architecture SYN_Behavioral of and2_264 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_263 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_263;

architecture SYN_Behavioral of and2_263 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_262 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_262;

architecture SYN_Behavioral of and2_262 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_261 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_261;

architecture SYN_Behavioral of and2_261 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_260 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_260;

architecture SYN_Behavioral of and2_260 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_259 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_259;

architecture SYN_Behavioral of and2_259 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_258 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_258;

architecture SYN_Behavioral of and2_258 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_257 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_257;

architecture SYN_Behavioral of and2_257 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_256 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_256;

architecture SYN_Behavioral of and2_256 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_255 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_255;

architecture SYN_Behavioral of and2_255 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_254 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_254;

architecture SYN_Behavioral of and2_254 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_253 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_253;

architecture SYN_Behavioral of and2_253 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_252 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_252;

architecture SYN_Behavioral of and2_252 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_251 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_251;

architecture SYN_Behavioral of and2_251 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_250 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_250;

architecture SYN_Behavioral of and2_250 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_249 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_249;

architecture SYN_Behavioral of and2_249 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_248 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_248;

architecture SYN_Behavioral of and2_248 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_247 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_247;

architecture SYN_Behavioral of and2_247 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_246 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_246;

architecture SYN_Behavioral of and2_246 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_245 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_245;

architecture SYN_Behavioral of and2_245 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_244 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_244;

architecture SYN_Behavioral of and2_244 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_243 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_243;

architecture SYN_Behavioral of and2_243 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_242 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_242;

architecture SYN_Behavioral of and2_242 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_241 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_241;

architecture SYN_Behavioral of and2_241 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_240 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_240;

architecture SYN_Behavioral of and2_240 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_239 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_239;

architecture SYN_Behavioral of and2_239 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_238 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_238;

architecture SYN_Behavioral of and2_238 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_237 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_237;

architecture SYN_Behavioral of and2_237 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_236 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_236;

architecture SYN_Behavioral of and2_236 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_235 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_235;

architecture SYN_Behavioral of and2_235 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_234 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_234;

architecture SYN_Behavioral of and2_234 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_233 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_233;

architecture SYN_Behavioral of and2_233 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_232 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_232;

architecture SYN_Behavioral of and2_232 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_231 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_231;

architecture SYN_Behavioral of and2_231 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_230 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_230;

architecture SYN_Behavioral of and2_230 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_229 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_229;

architecture SYN_Behavioral of and2_229 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_228 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_228;

architecture SYN_Behavioral of and2_228 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_227 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_227;

architecture SYN_Behavioral of and2_227 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_226 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_226;

architecture SYN_Behavioral of and2_226 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_225 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_225;

architecture SYN_Behavioral of and2_225 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_224 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_224;

architecture SYN_Behavioral of and2_224 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_223 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_223;

architecture SYN_Behavioral of and2_223 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_222 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_222;

architecture SYN_Behavioral of and2_222 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_221 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_221;

architecture SYN_Behavioral of and2_221 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_220 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_220;

architecture SYN_Behavioral of and2_220 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_219 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_219;

architecture SYN_Behavioral of and2_219 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_218 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_218;

architecture SYN_Behavioral of and2_218 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_217 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_217;

architecture SYN_Behavioral of and2_217 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_216 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_216;

architecture SYN_Behavioral of and2_216 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_215 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_215;

architecture SYN_Behavioral of and2_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_214 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_214;

architecture SYN_Behavioral of and2_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_213 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_213;

architecture SYN_Behavioral of and2_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_212 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_212;

architecture SYN_Behavioral of and2_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_211 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_211;

architecture SYN_Behavioral of and2_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_210 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_210;

architecture SYN_Behavioral of and2_210 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_209 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_209;

architecture SYN_Behavioral of and2_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_208 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_208;

architecture SYN_Behavioral of and2_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_207 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_207;

architecture SYN_Behavioral of and2_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_206 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_206;

architecture SYN_Behavioral of and2_206 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_205 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_205;

architecture SYN_Behavioral of and2_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_204 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_204;

architecture SYN_Behavioral of and2_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_203 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_203;

architecture SYN_Behavioral of and2_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_202 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_202;

architecture SYN_Behavioral of and2_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_201 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_201;

architecture SYN_Behavioral of and2_201 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_200 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_200;

architecture SYN_Behavioral of and2_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_199 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_199;

architecture SYN_Behavioral of and2_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_198 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_198;

architecture SYN_Behavioral of and2_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_197 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_197;

architecture SYN_Behavioral of and2_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_196 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_196;

architecture SYN_Behavioral of and2_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_195 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_195;

architecture SYN_Behavioral of and2_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_194 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_194;

architecture SYN_Behavioral of and2_194 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_193 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_193;

architecture SYN_Behavioral of and2_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_192 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_192;

architecture SYN_Behavioral of and2_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_191 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_191;

architecture SYN_Behavioral of and2_191 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_190 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_190;

architecture SYN_Behavioral of and2_190 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_189 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_189;

architecture SYN_Behavioral of and2_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_188 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_188;

architecture SYN_Behavioral of and2_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_187 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_187;

architecture SYN_Behavioral of and2_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_186 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_186;

architecture SYN_Behavioral of and2_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_185 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_185;

architecture SYN_Behavioral of and2_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_184 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_184;

architecture SYN_Behavioral of and2_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_183 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_183;

architecture SYN_Behavioral of and2_183 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_182 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_182;

architecture SYN_Behavioral of and2_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_181 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_181;

architecture SYN_Behavioral of and2_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_180 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_180;

architecture SYN_Behavioral of and2_180 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_179 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_179;

architecture SYN_Behavioral of and2_179 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_178 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_178;

architecture SYN_Behavioral of and2_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_177 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_177;

architecture SYN_Behavioral of and2_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_176 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_176;

architecture SYN_Behavioral of and2_176 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_175 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_175;

architecture SYN_Behavioral of and2_175 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_174 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_174;

architecture SYN_Behavioral of and2_174 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_173 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_173;

architecture SYN_Behavioral of and2_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_172 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_172;

architecture SYN_Behavioral of and2_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_171 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_171;

architecture SYN_Behavioral of and2_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_170 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_170;

architecture SYN_Behavioral of and2_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_169 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_169;

architecture SYN_Behavioral of and2_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_168 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_168;

architecture SYN_Behavioral of and2_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_167 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_167;

architecture SYN_Behavioral of and2_167 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_166 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_166;

architecture SYN_Behavioral of and2_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_165 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_165;

architecture SYN_Behavioral of and2_165 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_164 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_164;

architecture SYN_Behavioral of and2_164 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_163 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_163;

architecture SYN_Behavioral of and2_163 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_162 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_162;

architecture SYN_Behavioral of and2_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_161 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_161;

architecture SYN_Behavioral of and2_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_160 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_160;

architecture SYN_Behavioral of and2_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_159 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_159;

architecture SYN_Behavioral of and2_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_158 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_158;

architecture SYN_Behavioral of and2_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_157 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_157;

architecture SYN_Behavioral of and2_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_156 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_156;

architecture SYN_Behavioral of and2_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_155 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_155;

architecture SYN_Behavioral of and2_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_154 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_154;

architecture SYN_Behavioral of and2_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_153 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_153;

architecture SYN_Behavioral of and2_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_152 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_152;

architecture SYN_Behavioral of and2_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_151 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_151;

architecture SYN_Behavioral of and2_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_150 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_150;

architecture SYN_Behavioral of and2_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_149 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_149;

architecture SYN_Behavioral of and2_149 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_148 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_148;

architecture SYN_Behavioral of and2_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_147 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_147;

architecture SYN_Behavioral of and2_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_146 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_146;

architecture SYN_Behavioral of and2_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_145 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_145;

architecture SYN_Behavioral of and2_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_144 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_144;

architecture SYN_Behavioral of and2_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_143 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_143;

architecture SYN_Behavioral of and2_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_142 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_142;

architecture SYN_Behavioral of and2_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_141 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_141;

architecture SYN_Behavioral of and2_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_140 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_140;

architecture SYN_Behavioral of and2_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_139 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_139;

architecture SYN_Behavioral of and2_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_138 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_138;

architecture SYN_Behavioral of and2_138 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_137 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_137;

architecture SYN_Behavioral of and2_137 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_136 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_136;

architecture SYN_Behavioral of and2_136 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_135 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_135;

architecture SYN_Behavioral of and2_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_134 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_134;

architecture SYN_Behavioral of and2_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_133 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_133;

architecture SYN_Behavioral of and2_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_132 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_132;

architecture SYN_Behavioral of and2_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_131 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_131;

architecture SYN_Behavioral of and2_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_130 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_130;

architecture SYN_Behavioral of and2_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_129 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_129;

architecture SYN_Behavioral of and2_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_128 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_128;

architecture SYN_Behavioral of and2_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_127 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_127;

architecture SYN_Behavioral of and2_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_126 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_126;

architecture SYN_Behavioral of and2_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_125 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_125;

architecture SYN_Behavioral of and2_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_124 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_124;

architecture SYN_Behavioral of and2_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_123 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_123;

architecture SYN_Behavioral of and2_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_122 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_122;

architecture SYN_Behavioral of and2_122 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_121 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_121;

architecture SYN_Behavioral of and2_121 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_120 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_120;

architecture SYN_Behavioral of and2_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_119 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_119;

architecture SYN_Behavioral of and2_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_118 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_118;

architecture SYN_Behavioral of and2_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_117 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_117;

architecture SYN_Behavioral of and2_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_116 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_116;

architecture SYN_Behavioral of and2_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_115 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_115;

architecture SYN_Behavioral of and2_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_114 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_114;

architecture SYN_Behavioral of and2_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_113 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_113;

architecture SYN_Behavioral of and2_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_112 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_112;

architecture SYN_Behavioral of and2_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_111 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_111;

architecture SYN_Behavioral of and2_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_110 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_110;

architecture SYN_Behavioral of and2_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_109 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_109;

architecture SYN_Behavioral of and2_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_108 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_108;

architecture SYN_Behavioral of and2_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_107 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_107;

architecture SYN_Behavioral of and2_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_106 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_106;

architecture SYN_Behavioral of and2_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_105 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_105;

architecture SYN_Behavioral of and2_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_104 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_104;

architecture SYN_Behavioral of and2_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_103 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_103;

architecture SYN_Behavioral of and2_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_102 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_102;

architecture SYN_Behavioral of and2_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_101 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_101;

architecture SYN_Behavioral of and2_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_100 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_100;

architecture SYN_Behavioral of and2_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_99 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_99;

architecture SYN_Behavioral of and2_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_98 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_98;

architecture SYN_Behavioral of and2_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_97 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_97;

architecture SYN_Behavioral of and2_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_96 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_96;

architecture SYN_Behavioral of and2_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_95 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_95;

architecture SYN_Behavioral of and2_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_94 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_94;

architecture SYN_Behavioral of and2_94 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_93 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_93;

architecture SYN_Behavioral of and2_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_92 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_92;

architecture SYN_Behavioral of and2_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_91 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_91;

architecture SYN_Behavioral of and2_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_90 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_90;

architecture SYN_Behavioral of and2_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_89 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_89;

architecture SYN_Behavioral of and2_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_88 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_88;

architecture SYN_Behavioral of and2_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_87 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_87;

architecture SYN_Behavioral of and2_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_86 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_86;

architecture SYN_Behavioral of and2_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_85 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_85;

architecture SYN_Behavioral of and2_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_84 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_84;

architecture SYN_Behavioral of and2_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_83 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_83;

architecture SYN_Behavioral of and2_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_82 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_82;

architecture SYN_Behavioral of and2_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_81 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_81;

architecture SYN_Behavioral of and2_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_80 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_80;

architecture SYN_Behavioral of and2_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_79 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_79;

architecture SYN_Behavioral of and2_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_78 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_78;

architecture SYN_Behavioral of and2_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_77 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_77;

architecture SYN_Behavioral of and2_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_76 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_76;

architecture SYN_Behavioral of and2_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_75 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_75;

architecture SYN_Behavioral of and2_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_74 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_74;

architecture SYN_Behavioral of and2_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_73 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_73;

architecture SYN_Behavioral of and2_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_72 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_72;

architecture SYN_Behavioral of and2_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_71 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_71;

architecture SYN_Behavioral of and2_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_70 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_70;

architecture SYN_Behavioral of and2_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_69 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_69;

architecture SYN_Behavioral of and2_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_68 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_68;

architecture SYN_Behavioral of and2_68 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_67 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_67;

architecture SYN_Behavioral of and2_67 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_66 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_66;

architecture SYN_Behavioral of and2_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_65 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_65;

architecture SYN_Behavioral of and2_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_64 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_64;

architecture SYN_Behavioral of and2_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_63 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_63;

architecture SYN_Behavioral of and2_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_62 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_62;

architecture SYN_Behavioral of and2_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_61 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_61;

architecture SYN_Behavioral of and2_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_60 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_60;

architecture SYN_Behavioral of and2_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_59 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_59;

architecture SYN_Behavioral of and2_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_58 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_58;

architecture SYN_Behavioral of and2_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_57 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_57;

architecture SYN_Behavioral of and2_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_56 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_56;

architecture SYN_Behavioral of and2_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_55 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_55;

architecture SYN_Behavioral of and2_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_54 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_54;

architecture SYN_Behavioral of and2_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_53 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_53;

architecture SYN_Behavioral of and2_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_52 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_52;

architecture SYN_Behavioral of and2_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_51 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_51;

architecture SYN_Behavioral of and2_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_50 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_50;

architecture SYN_Behavioral of and2_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_49 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_49;

architecture SYN_Behavioral of and2_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_48 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_48;

architecture SYN_Behavioral of and2_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_47 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_47;

architecture SYN_Behavioral of and2_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_46 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_46;

architecture SYN_Behavioral of and2_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_45 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_45;

architecture SYN_Behavioral of and2_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_44 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_44;

architecture SYN_Behavioral of and2_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_43 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_43;

architecture SYN_Behavioral of and2_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_42 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_42;

architecture SYN_Behavioral of and2_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_41 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_41;

architecture SYN_Behavioral of and2_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_40 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_40;

architecture SYN_Behavioral of and2_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_39 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_39;

architecture SYN_Behavioral of and2_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_38 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_38;

architecture SYN_Behavioral of and2_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_37 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_37;

architecture SYN_Behavioral of and2_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_36 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_36;

architecture SYN_Behavioral of and2_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_35 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_35;

architecture SYN_Behavioral of and2_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_34 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_34;

architecture SYN_Behavioral of and2_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_33 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_33;

architecture SYN_Behavioral of and2_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_32 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_32;

architecture SYN_Behavioral of and2_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_31 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_31;

architecture SYN_Behavioral of and2_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_30 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_30;

architecture SYN_Behavioral of and2_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_29 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_29;

architecture SYN_Behavioral of and2_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_28 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_28;

architecture SYN_Behavioral of and2_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_27 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_27;

architecture SYN_Behavioral of and2_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_26 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_26;

architecture SYN_Behavioral of and2_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_25 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_25;

architecture SYN_Behavioral of and2_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_24 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_24;

architecture SYN_Behavioral of and2_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_23 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_23;

architecture SYN_Behavioral of and2_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_22 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_22;

architecture SYN_Behavioral of and2_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_21 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_21;

architecture SYN_Behavioral of and2_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_20 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_20;

architecture SYN_Behavioral of and2_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_19 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_19;

architecture SYN_Behavioral of and2_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_18 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_18;

architecture SYN_Behavioral of and2_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_17 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_17;

architecture SYN_Behavioral of and2_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_16 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_16;

architecture SYN_Behavioral of and2_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_15 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_15;

architecture SYN_Behavioral of and2_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_14 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_14;

architecture SYN_Behavioral of and2_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_13 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_13;

architecture SYN_Behavioral of and2_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_12 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_12;

architecture SYN_Behavioral of and2_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_11 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_11;

architecture SYN_Behavioral of and2_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_10 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_10;

architecture SYN_Behavioral of and2_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_9 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_9;

architecture SYN_Behavioral of and2_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_8 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_8;

architecture SYN_Behavioral of and2_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_7 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_7;

architecture SYN_Behavioral of and2_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_6 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_6;

architecture SYN_Behavioral of and2_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_5 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_5;

architecture SYN_Behavioral of and2_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_4 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_4;

architecture SYN_Behavioral of and2_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_3 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_3;

architecture SYN_Behavioral of and2_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_2 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_2;

architecture SYN_Behavioral of and2_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_1 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_1;

architecture SYN_Behavioral of and2_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_63 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_63;

architecture SYN_full_adder_arc of full_adder_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_62 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_62;

architecture SYN_full_adder_arc of full_adder_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_61 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_61;

architecture SYN_full_adder_arc of full_adder_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_60 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_60;

architecture SYN_full_adder_arc of full_adder_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_59 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_59;

architecture SYN_full_adder_arc of full_adder_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_58 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_58;

architecture SYN_full_adder_arc of full_adder_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_57 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_57;

architecture SYN_full_adder_arc of full_adder_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_56 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_56;

architecture SYN_full_adder_arc of full_adder_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_55 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_55;

architecture SYN_full_adder_arc of full_adder_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_54 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_54;

architecture SYN_full_adder_arc of full_adder_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_53 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_53;

architecture SYN_full_adder_arc of full_adder_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_52 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_52;

architecture SYN_full_adder_arc of full_adder_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_51 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_51;

architecture SYN_full_adder_arc of full_adder_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_50 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_50;

architecture SYN_full_adder_arc of full_adder_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_49 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_49;

architecture SYN_full_adder_arc of full_adder_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_48 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_48;

architecture SYN_full_adder_arc of full_adder_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_47 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_47;

architecture SYN_full_adder_arc of full_adder_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_46 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_46;

architecture SYN_full_adder_arc of full_adder_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_45 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_45;

architecture SYN_full_adder_arc of full_adder_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_44 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_44;

architecture SYN_full_adder_arc of full_adder_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_43 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_43;

architecture SYN_full_adder_arc of full_adder_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_42 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_42;

architecture SYN_full_adder_arc of full_adder_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_41 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_41;

architecture SYN_full_adder_arc of full_adder_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_40 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_40;

architecture SYN_full_adder_arc of full_adder_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_39 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_39;

architecture SYN_full_adder_arc of full_adder_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_38 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_38;

architecture SYN_full_adder_arc of full_adder_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_37 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_37;

architecture SYN_full_adder_arc of full_adder_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_36 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_36;

architecture SYN_full_adder_arc of full_adder_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_35 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_35;

architecture SYN_full_adder_arc of full_adder_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_34 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_34;

architecture SYN_full_adder_arc of full_adder_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_33 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_33;

architecture SYN_full_adder_arc of full_adder_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_32 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_32;

architecture SYN_full_adder_arc of full_adder_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_31 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_31;

architecture SYN_full_adder_arc of full_adder_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_30 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_30;

architecture SYN_full_adder_arc of full_adder_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_29 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_29;

architecture SYN_full_adder_arc of full_adder_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_28 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_28;

architecture SYN_full_adder_arc of full_adder_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_27 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_27;

architecture SYN_full_adder_arc of full_adder_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_26 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_26;

architecture SYN_full_adder_arc of full_adder_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_25 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_25;

architecture SYN_full_adder_arc of full_adder_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_24 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_24;

architecture SYN_full_adder_arc of full_adder_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_23 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_23;

architecture SYN_full_adder_arc of full_adder_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_22 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_22;

architecture SYN_full_adder_arc of full_adder_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_21 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_21;

architecture SYN_full_adder_arc of full_adder_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_20 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_20;

architecture SYN_full_adder_arc of full_adder_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_19 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_19;

architecture SYN_full_adder_arc of full_adder_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_18 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_18;

architecture SYN_full_adder_arc of full_adder_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_17 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_17;

architecture SYN_full_adder_arc of full_adder_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_16 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_16;

architecture SYN_full_adder_arc of full_adder_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_15 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_15;

architecture SYN_full_adder_arc of full_adder_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_14 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_14;

architecture SYN_full_adder_arc of full_adder_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_13 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_13;

architecture SYN_full_adder_arc of full_adder_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_12 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_12;

architecture SYN_full_adder_arc of full_adder_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_11 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_11;

architecture SYN_full_adder_arc of full_adder_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_10 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_10;

architecture SYN_full_adder_arc of full_adder_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_9 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_9;

architecture SYN_full_adder_arc of full_adder_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_8 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_8;

architecture SYN_full_adder_arc of full_adder_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_7 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_7;

architecture SYN_full_adder_arc of full_adder_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_6 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_6;

architecture SYN_full_adder_arc of full_adder_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_5 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_5;

architecture SYN_full_adder_arc of full_adder_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_4 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_4;

architecture SYN_full_adder_arc of full_adder_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_3 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_3;

architecture SYN_full_adder_arc of full_adder_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_2 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_2;

architecture SYN_full_adder_arc of full_adder_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_1 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_1;

architecture SYN_full_adder_arc of full_adder_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_216 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_216;

architecture SYN_Structural of fa_216 is

   component or2_216
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_437
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_438
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_437
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_438
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_438 port map( a => a, b => b, o => s1);
   xor_2 : xor2_437 port map( a => s1, b => ci, o => s);
   and_1 : and2_438 port map( a => a, b => b, o => s2);
   and_2 : and2_437 port map( a => s1, b => ci, o => s3);
   or_1 : or2_216 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_215 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_215;

architecture SYN_Structural of fa_215 is

   component or2_215
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_435
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_436
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_435
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_436
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_436 port map( a => a, b => b, o => s1);
   xor_2 : xor2_435 port map( a => s1, b => ci, o => s);
   and_1 : and2_436 port map( a => a, b => b, o => s2);
   and_2 : and2_435 port map( a => s1, b => ci, o => s3);
   or_1 : or2_215 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_214 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_214;

architecture SYN_Structural of fa_214 is

   component or2_214
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_433
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_434
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_433
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_434
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_434 port map( a => a, b => b, o => s1);
   xor_2 : xor2_433 port map( a => s1, b => ci, o => s);
   and_1 : and2_434 port map( a => a, b => b, o => s2);
   and_2 : and2_433 port map( a => s1, b => ci, o => s3);
   or_1 : or2_214 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_213 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_213;

architecture SYN_Structural of fa_213 is

   component or2_213
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_431
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_432
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_431
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_432
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_432 port map( a => a, b => b, o => s1);
   xor_2 : xor2_431 port map( a => s1, b => ci, o => s);
   and_1 : and2_432 port map( a => a, b => b, o => s2);
   and_2 : and2_431 port map( a => s1, b => ci, o => s3);
   or_1 : or2_213 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_212 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_212;

architecture SYN_Structural of fa_212 is

   component or2_212
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_429
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_430
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_429
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_430
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_430 port map( a => a, b => b, o => s1);
   xor_2 : xor2_429 port map( a => s1, b => ci, o => s);
   and_1 : and2_430 port map( a => a, b => b, o => s2);
   and_2 : and2_429 port map( a => s1, b => ci, o => s3);
   or_1 : or2_212 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_211 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_211;

architecture SYN_Structural of fa_211 is

   component or2_211
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_427
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_428
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_427
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_428
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_428 port map( a => a, b => b, o => s1);
   xor_2 : xor2_427 port map( a => s1, b => ci, o => s);
   and_1 : and2_428 port map( a => a, b => b, o => s2);
   and_2 : and2_427 port map( a => s1, b => ci, o => s3);
   or_1 : or2_211 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_210 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_210;

architecture SYN_Structural of fa_210 is

   component or2_210
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_425
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_426
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_425
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_426
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_426 port map( a => a, b => b, o => s1);
   xor_2 : xor2_425 port map( a => s1, b => ci, o => s);
   and_1 : and2_426 port map( a => a, b => b, o => s2);
   and_2 : and2_425 port map( a => s1, b => ci, o => s3);
   or_1 : or2_210 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_209 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_209;

architecture SYN_Structural of fa_209 is

   component or2_209
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_423
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_424
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_423
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_424
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_424 port map( a => a, b => b, o => s1);
   xor_2 : xor2_423 port map( a => s1, b => ci, o => s);
   and_1 : and2_424 port map( a => a, b => b, o => s2);
   and_2 : and2_423 port map( a => s1, b => ci, o => s3);
   or_1 : or2_209 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_208 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_208;

architecture SYN_Structural of fa_208 is

   component or2_208
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_421
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_422
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_421
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_422
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_422 port map( a => a, b => b, o => s1);
   xor_2 : xor2_421 port map( a => s1, b => ci, o => s);
   and_1 : and2_422 port map( a => a, b => b, o => s2);
   and_2 : and2_421 port map( a => s1, b => ci, o => s3);
   or_1 : or2_208 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_207 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_207;

architecture SYN_Structural of fa_207 is

   component or2_207
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_419
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_420
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_419
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_420
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_420 port map( a => a, b => b, o => s1);
   xor_2 : xor2_419 port map( a => s1, b => ci, o => s);
   and_1 : and2_420 port map( a => a, b => b, o => s2);
   and_2 : and2_419 port map( a => s1, b => ci, o => s3);
   or_1 : or2_207 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_206 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_206;

architecture SYN_Structural of fa_206 is

   component or2_206
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_417
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_418
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_417
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_418
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_418 port map( a => a, b => b, o => s1);
   xor_2 : xor2_417 port map( a => s1, b => ci, o => s);
   and_1 : and2_418 port map( a => a, b => b, o => s2);
   and_2 : and2_417 port map( a => s1, b => ci, o => s3);
   or_1 : or2_206 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_205 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_205;

architecture SYN_Structural of fa_205 is

   component or2_205
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_415
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_416
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_415
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_416
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_416 port map( a => a, b => b, o => s1);
   xor_2 : xor2_415 port map( a => s1, b => ci, o => s);
   and_1 : and2_416 port map( a => a, b => b, o => s2);
   and_2 : and2_415 port map( a => s1, b => ci, o => s3);
   or_1 : or2_205 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_204 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_204;

architecture SYN_Structural of fa_204 is

   component or2_204
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_413
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_414
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_413
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_414
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_414 port map( a => a, b => b, o => s1);
   xor_2 : xor2_413 port map( a => s1, b => ci, o => s);
   and_1 : and2_414 port map( a => a, b => b, o => s2);
   and_2 : and2_413 port map( a => s1, b => ci, o => s3);
   or_1 : or2_204 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_203 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_203;

architecture SYN_Structural of fa_203 is

   component or2_203
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_411
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_412
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_411
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_412
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_412 port map( a => a, b => b, o => s1);
   xor_2 : xor2_411 port map( a => s1, b => ci, o => s);
   and_1 : and2_412 port map( a => a, b => b, o => s2);
   and_2 : and2_411 port map( a => s1, b => ci, o => s3);
   or_1 : or2_203 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_202 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_202;

architecture SYN_Structural of fa_202 is

   component or2_202
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_409
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_410
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_409
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_410
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_410 port map( a => a, b => b, o => s1);
   xor_2 : xor2_409 port map( a => s1, b => ci, o => s);
   and_1 : and2_410 port map( a => a, b => b, o => s2);
   and_2 : and2_409 port map( a => s1, b => ci, o => s3);
   or_1 : or2_202 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_201 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_201;

architecture SYN_Structural of fa_201 is

   component or2_201
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_407
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_408
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_407
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_408
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_408 port map( a => a, b => b, o => s1);
   xor_2 : xor2_407 port map( a => s1, b => ci, o => s);
   and_1 : and2_408 port map( a => a, b => b, o => s2);
   and_2 : and2_407 port map( a => s1, b => ci, o => s3);
   or_1 : or2_201 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_200 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_200;

architecture SYN_Structural of fa_200 is

   component or2_200
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_405
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_406
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_405
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_406
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_406 port map( a => a, b => b, o => s1);
   xor_2 : xor2_405 port map( a => s1, b => ci, o => s);
   and_1 : and2_406 port map( a => a, b => b, o => s2);
   and_2 : and2_405 port map( a => s1, b => ci, o => s3);
   or_1 : or2_200 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_199 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_199;

architecture SYN_Structural of fa_199 is

   component or2_199
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_403
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_404
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_403
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_404
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_404 port map( a => a, b => b, o => s1);
   xor_2 : xor2_403 port map( a => s1, b => ci, o => s);
   and_1 : and2_404 port map( a => a, b => b, o => s2);
   and_2 : and2_403 port map( a => s1, b => ci, o => s3);
   or_1 : or2_199 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_198 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_198;

architecture SYN_Structural of fa_198 is

   component or2_198
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_401
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_402
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_401
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_402
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_402 port map( a => a, b => b, o => s1);
   xor_2 : xor2_401 port map( a => s1, b => ci, o => s);
   and_1 : and2_402 port map( a => a, b => b, o => s2);
   and_2 : and2_401 port map( a => s1, b => ci, o => s3);
   or_1 : or2_198 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_197 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_197;

architecture SYN_Structural of fa_197 is

   component or2_197
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_399
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_400
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_399
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_400
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_400 port map( a => a, b => b, o => s1);
   xor_2 : xor2_399 port map( a => s1, b => ci, o => s);
   and_1 : and2_400 port map( a => a, b => b, o => s2);
   and_2 : and2_399 port map( a => s1, b => ci, o => s3);
   or_1 : or2_197 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_196 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_196;

architecture SYN_Structural of fa_196 is

   component or2_196
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_397
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_398
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_397
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_398
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_398 port map( a => a, b => b, o => s1);
   xor_2 : xor2_397 port map( a => s1, b => ci, o => s);
   and_1 : and2_398 port map( a => a, b => b, o => s2);
   and_2 : and2_397 port map( a => s1, b => ci, o => s3);
   or_1 : or2_196 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_195 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_195;

architecture SYN_Structural of fa_195 is

   component or2_195
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_395
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_396
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_395
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_396
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_396 port map( a => a, b => b, o => s1);
   xor_2 : xor2_395 port map( a => s1, b => ci, o => s);
   and_1 : and2_396 port map( a => a, b => b, o => s2);
   and_2 : and2_395 port map( a => s1, b => ci, o => s3);
   or_1 : or2_195 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_194 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_194;

architecture SYN_Structural of fa_194 is

   component or2_194
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_393
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_394
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_393
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_394
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_394 port map( a => a, b => b, o => s1);
   xor_2 : xor2_393 port map( a => s1, b => ci, o => s);
   and_1 : and2_394 port map( a => a, b => b, o => s2);
   and_2 : and2_393 port map( a => s1, b => ci, o => s3);
   or_1 : or2_194 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_193 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_193;

architecture SYN_Structural of fa_193 is

   component or2_193
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_391
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_392
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_391
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_392
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_392 port map( a => a, b => b, o => s1);
   xor_2 : xor2_391 port map( a => s1, b => ci, o => s);
   and_1 : and2_392 port map( a => a, b => b, o => s2);
   and_2 : and2_391 port map( a => s1, b => ci, o => s3);
   or_1 : or2_193 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_192 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_192;

architecture SYN_Structural of fa_192 is

   component or2_192
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_389
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_390
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_389
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_390
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_390 port map( a => a, b => b, o => s1);
   xor_2 : xor2_389 port map( a => s1, b => ci, o => s);
   and_1 : and2_390 port map( a => a, b => b, o => s2);
   and_2 : and2_389 port map( a => s1, b => ci, o => s3);
   or_1 : or2_192 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_191 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_191;

architecture SYN_Structural of fa_191 is

   component or2_191
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_387
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_388
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_387
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_388
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_388 port map( a => a, b => b, o => s1);
   xor_2 : xor2_387 port map( a => s1, b => ci, o => s);
   and_1 : and2_388 port map( a => a, b => b, o => s2);
   and_2 : and2_387 port map( a => s1, b => ci, o => s3);
   or_1 : or2_191 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_190 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_190;

architecture SYN_Structural of fa_190 is

   component or2_190
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_385
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_386
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_385
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_386
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_386 port map( a => a, b => b, o => s1);
   xor_2 : xor2_385 port map( a => s1, b => ci, o => s);
   and_1 : and2_386 port map( a => a, b => b, o => s2);
   and_2 : and2_385 port map( a => s1, b => ci, o => s3);
   or_1 : or2_190 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_189 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_189;

architecture SYN_Structural of fa_189 is

   component or2_189
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_383
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_384
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_383
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_384
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_384 port map( a => a, b => b, o => s1);
   xor_2 : xor2_383 port map( a => s1, b => ci, o => s);
   and_1 : and2_384 port map( a => a, b => b, o => s2);
   and_2 : and2_383 port map( a => s1, b => ci, o => s3);
   or_1 : or2_189 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_188 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_188;

architecture SYN_Structural of fa_188 is

   component or2_188
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_381
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_382
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_381
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_382
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_382 port map( a => a, b => b, o => s1);
   xor_2 : xor2_381 port map( a => s1, b => ci, o => s);
   and_1 : and2_382 port map( a => a, b => b, o => s2);
   and_2 : and2_381 port map( a => s1, b => ci, o => s3);
   or_1 : or2_188 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_187 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_187;

architecture SYN_Structural of fa_187 is

   component or2_187
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_379
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_380
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_379
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_380
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_380 port map( a => a, b => b, o => s1);
   xor_2 : xor2_379 port map( a => s1, b => ci, o => s);
   and_1 : and2_380 port map( a => a, b => b, o => s2);
   and_2 : and2_379 port map( a => s1, b => ci, o => s3);
   or_1 : or2_187 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_186 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_186;

architecture SYN_Structural of fa_186 is

   component or2_186
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_376
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_377
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_376
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_377
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_377 port map( a => a, b => b, o => s1);
   xor_2 : xor2_376 port map( a => s1, b => ci, o => s);
   and_1 : and2_377 port map( a => a, b => b, o => s2);
   and_2 : and2_376 port map( a => s1, b => ci, o => s3);
   or_1 : or2_186 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_185 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_185;

architecture SYN_Structural of fa_185 is

   component or2_185
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_374
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_375
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_374
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_375
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_375 port map( a => a, b => b, o => s1);
   xor_2 : xor2_374 port map( a => s1, b => ci, o => s);
   and_1 : and2_375 port map( a => a, b => b, o => s2);
   and_2 : and2_374 port map( a => s1, b => ci, o => s3);
   or_1 : or2_185 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_184 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_184;

architecture SYN_Structural of fa_184 is

   component or2_184
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_372
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_373
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_372
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_373
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_373 port map( a => a, b => b, o => s1);
   xor_2 : xor2_372 port map( a => s1, b => ci, o => s);
   and_1 : and2_373 port map( a => a, b => b, o => s2);
   and_2 : and2_372 port map( a => s1, b => ci, o => s3);
   or_1 : or2_184 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_183 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_183;

architecture SYN_Structural of fa_183 is

   component or2_183
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_370
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_371
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_370
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_371
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_371 port map( a => a, b => b, o => s1);
   xor_2 : xor2_370 port map( a => s1, b => ci, o => s);
   and_1 : and2_371 port map( a => a, b => b, o => s2);
   and_2 : and2_370 port map( a => s1, b => ci, o => s3);
   or_1 : or2_183 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_182 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_182;

architecture SYN_Structural of fa_182 is

   component or2_182
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_368
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_369
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_368
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_369
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_369 port map( a => a, b => b, o => s1);
   xor_2 : xor2_368 port map( a => s1, b => ci, o => s);
   and_1 : and2_369 port map( a => a, b => b, o => s2);
   and_2 : and2_368 port map( a => s1, b => ci, o => s3);
   or_1 : or2_182 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_181 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_181;

architecture SYN_Structural of fa_181 is

   component or2_181
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_366
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_367
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_366
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_367
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_367 port map( a => a, b => b, o => s1);
   xor_2 : xor2_366 port map( a => s1, b => ci, o => s);
   and_1 : and2_367 port map( a => a, b => b, o => s2);
   and_2 : and2_366 port map( a => s1, b => ci, o => s3);
   or_1 : or2_181 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_180 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_180;

architecture SYN_Structural of fa_180 is

   component or2_180
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_364
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_365
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_364
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_365
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_365 port map( a => a, b => b, o => s1);
   xor_2 : xor2_364 port map( a => s1, b => ci, o => s);
   and_1 : and2_365 port map( a => a, b => b, o => s2);
   and_2 : and2_364 port map( a => s1, b => ci, o => s3);
   or_1 : or2_180 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_179 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_179;

architecture SYN_Structural of fa_179 is

   component or2_179
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_362
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_363
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_362
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_363
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_363 port map( a => a, b => b, o => s1);
   xor_2 : xor2_362 port map( a => s1, b => ci, o => s);
   and_1 : and2_363 port map( a => a, b => b, o => s2);
   and_2 : and2_362 port map( a => s1, b => ci, o => s3);
   or_1 : or2_179 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_178 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_178;

architecture SYN_Structural of fa_178 is

   component or2_178
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_360
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_361
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_360
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_361
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_361 port map( a => a, b => b, o => s1);
   xor_2 : xor2_360 port map( a => s1, b => ci, o => s);
   and_1 : and2_361 port map( a => a, b => b, o => s2);
   and_2 : and2_360 port map( a => s1, b => ci, o => s3);
   or_1 : or2_178 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_177 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_177;

architecture SYN_Structural of fa_177 is

   component or2_177
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_358
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_359
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_358
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_359
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_359 port map( a => a, b => b, o => s1);
   xor_2 : xor2_358 port map( a => s1, b => ci, o => s);
   and_1 : and2_359 port map( a => a, b => b, o => s2);
   and_2 : and2_358 port map( a => s1, b => ci, o => s3);
   or_1 : or2_177 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_176 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_176;

architecture SYN_Structural of fa_176 is

   component or2_176
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_356
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_357
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_356
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_357
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_357 port map( a => a, b => b, o => s1);
   xor_2 : xor2_356 port map( a => s1, b => ci, o => s);
   and_1 : and2_357 port map( a => a, b => b, o => s2);
   and_2 : and2_356 port map( a => s1, b => ci, o => s3);
   or_1 : or2_176 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_175 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_175;

architecture SYN_Structural of fa_175 is

   component or2_175
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_354
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_355
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_354
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_355
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_355 port map( a => a, b => b, o => s1);
   xor_2 : xor2_354 port map( a => s1, b => ci, o => s);
   and_1 : and2_355 port map( a => a, b => b, o => s2);
   and_2 : and2_354 port map( a => s1, b => ci, o => s3);
   or_1 : or2_175 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_174 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_174;

architecture SYN_Structural of fa_174 is

   component or2_174
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_352
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_353
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_352
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_353
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_353 port map( a => a, b => b, o => s1);
   xor_2 : xor2_352 port map( a => s1, b => ci, o => s);
   and_1 : and2_353 port map( a => a, b => b, o => s2);
   and_2 : and2_352 port map( a => s1, b => ci, o => s3);
   or_1 : or2_174 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_173 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_173;

architecture SYN_Structural of fa_173 is

   component or2_173
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_350
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_351
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_350
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_351
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_351 port map( a => a, b => b, o => s1);
   xor_2 : xor2_350 port map( a => s1, b => ci, o => s);
   and_1 : and2_351 port map( a => a, b => b, o => s2);
   and_2 : and2_350 port map( a => s1, b => ci, o => s3);
   or_1 : or2_173 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_172 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_172;

architecture SYN_Structural of fa_172 is

   component or2_172
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_348
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_349
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_348
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_349
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_349 port map( a => a, b => b, o => s1);
   xor_2 : xor2_348 port map( a => s1, b => ci, o => s);
   and_1 : and2_349 port map( a => a, b => b, o => s2);
   and_2 : and2_348 port map( a => s1, b => ci, o => s3);
   or_1 : or2_172 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_171 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_171;

architecture SYN_Structural of fa_171 is

   component or2_171
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_346
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_347
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_346
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_347
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_347 port map( a => a, b => b, o => s1);
   xor_2 : xor2_346 port map( a => s1, b => ci, o => s);
   and_1 : and2_347 port map( a => a, b => b, o => s2);
   and_2 : and2_346 port map( a => s1, b => ci, o => s3);
   or_1 : or2_171 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_170 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_170;

architecture SYN_Structural of fa_170 is

   component or2_170
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_344
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_345
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_344
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_345
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_345 port map( a => a, b => b, o => s1);
   xor_2 : xor2_344 port map( a => s1, b => ci, o => s);
   and_1 : and2_345 port map( a => a, b => b, o => s2);
   and_2 : and2_344 port map( a => s1, b => ci, o => s3);
   or_1 : or2_170 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_169 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_169;

architecture SYN_Structural of fa_169 is

   component or2_169
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_342
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_343
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_342
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_343
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_343 port map( a => a, b => b, o => s1);
   xor_2 : xor2_342 port map( a => s1, b => ci, o => s);
   and_1 : and2_343 port map( a => a, b => b, o => s2);
   and_2 : and2_342 port map( a => s1, b => ci, o => s3);
   or_1 : or2_169 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_168 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_168;

architecture SYN_Structural of fa_168 is

   component or2_168
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_340
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_341
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_340
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_341
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_341 port map( a => a, b => b, o => s1);
   xor_2 : xor2_340 port map( a => s1, b => ci, o => s);
   and_1 : and2_341 port map( a => a, b => b, o => s2);
   and_2 : and2_340 port map( a => s1, b => ci, o => s3);
   or_1 : or2_168 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_167 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_167;

architecture SYN_Structural of fa_167 is

   component or2_167
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_338
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_339
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_338
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_339
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_339 port map( a => a, b => b, o => s1);
   xor_2 : xor2_338 port map( a => s1, b => ci, o => s);
   and_1 : and2_339 port map( a => a, b => b, o => s2);
   and_2 : and2_338 port map( a => s1, b => ci, o => s3);
   or_1 : or2_167 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_166 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_166;

architecture SYN_Structural of fa_166 is

   component or2_166
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_336
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_337
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_336
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_337
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_337 port map( a => a, b => b, o => s1);
   xor_2 : xor2_336 port map( a => s1, b => ci, o => s);
   and_1 : and2_337 port map( a => a, b => b, o => s2);
   and_2 : and2_336 port map( a => s1, b => ci, o => s3);
   or_1 : or2_166 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_165 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_165;

architecture SYN_Structural of fa_165 is

   component or2_165
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_334
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_335
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_334
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_335
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_335 port map( a => a, b => b, o => s1);
   xor_2 : xor2_334 port map( a => s1, b => ci, o => s);
   and_1 : and2_335 port map( a => a, b => b, o => s2);
   and_2 : and2_334 port map( a => s1, b => ci, o => s3);
   or_1 : or2_165 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_164 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_164;

architecture SYN_Structural of fa_164 is

   component or2_164
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_332
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_333
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_332
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_333
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_333 port map( a => a, b => b, o => s1);
   xor_2 : xor2_332 port map( a => s1, b => ci, o => s);
   and_1 : and2_333 port map( a => a, b => b, o => s2);
   and_2 : and2_332 port map( a => s1, b => ci, o => s3);
   or_1 : or2_164 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_163 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_163;

architecture SYN_Structural of fa_163 is

   component or2_163
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_330
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_331
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_330
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_331
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_331 port map( a => a, b => b, o => s1);
   xor_2 : xor2_330 port map( a => s1, b => ci, o => s);
   and_1 : and2_331 port map( a => a, b => b, o => s2);
   and_2 : and2_330 port map( a => s1, b => ci, o => s3);
   or_1 : or2_163 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_162 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_162;

architecture SYN_Structural of fa_162 is

   component or2_162
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_328
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_329
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_328
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_329
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_329 port map( a => a, b => b, o => s1);
   xor_2 : xor2_328 port map( a => s1, b => ci, o => s);
   and_1 : and2_329 port map( a => a, b => b, o => s2);
   and_2 : and2_328 port map( a => s1, b => ci, o => s3);
   or_1 : or2_162 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_161 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_161;

architecture SYN_Structural of fa_161 is

   component or2_161
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_326
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_327
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_326
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_327
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_327 port map( a => a, b => b, o => s1);
   xor_2 : xor2_326 port map( a => s1, b => ci, o => s);
   and_1 : and2_327 port map( a => a, b => b, o => s2);
   and_2 : and2_326 port map( a => s1, b => ci, o => s3);
   or_1 : or2_161 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_160 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_160;

architecture SYN_Structural of fa_160 is

   component or2_160
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_324
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_325
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_324
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_325
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_325 port map( a => a, b => b, o => s1);
   xor_2 : xor2_324 port map( a => s1, b => ci, o => s);
   and_1 : and2_325 port map( a => a, b => b, o => s2);
   and_2 : and2_324 port map( a => s1, b => ci, o => s3);
   or_1 : or2_160 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_159 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_159;

architecture SYN_Structural of fa_159 is

   component or2_159
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_322
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_323
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_322
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_323
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_323 port map( a => a, b => b, o => s1);
   xor_2 : xor2_322 port map( a => s1, b => ci, o => s);
   and_1 : and2_323 port map( a => a, b => b, o => s2);
   and_2 : and2_322 port map( a => s1, b => ci, o => s3);
   or_1 : or2_159 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_158 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_158;

architecture SYN_Structural of fa_158 is

   component or2_158
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_320
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_321
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_320
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_321
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_321 port map( a => a, b => b, o => s1);
   xor_2 : xor2_320 port map( a => s1, b => ci, o => s);
   and_1 : and2_321 port map( a => a, b => b, o => s2);
   and_2 : and2_320 port map( a => s1, b => ci, o => s3);
   or_1 : or2_158 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_157 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_157;

architecture SYN_Structural of fa_157 is

   component or2_157
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_318
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_319
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_318
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_319
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_319 port map( a => a, b => b, o => s1);
   xor_2 : xor2_318 port map( a => s1, b => ci, o => s);
   and_1 : and2_319 port map( a => a, b => b, o => s2);
   and_2 : and2_318 port map( a => s1, b => ci, o => s3);
   or_1 : or2_157 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_156 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_156;

architecture SYN_Structural of fa_156 is

   component or2_156
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_316
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_317
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_316
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_317
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_317 port map( a => a, b => b, o => s1);
   xor_2 : xor2_316 port map( a => s1, b => ci, o => s);
   and_1 : and2_317 port map( a => a, b => b, o => s2);
   and_2 : and2_316 port map( a => s1, b => ci, o => s3);
   or_1 : or2_156 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_155 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_155;

architecture SYN_Structural of fa_155 is

   component or2_155
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_313
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_314
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_313
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_314
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_314 port map( a => a, b => b, o => s1);
   xor_2 : xor2_313 port map( a => s1, b => ci, o => s);
   and_1 : and2_314 port map( a => a, b => b, o => s2);
   and_2 : and2_313 port map( a => s1, b => ci, o => s3);
   or_1 : or2_155 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_154 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_154;

architecture SYN_Structural of fa_154 is

   component or2_154
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_311
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_312
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_311
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_312
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_312 port map( a => a, b => b, o => s1);
   xor_2 : xor2_311 port map( a => s1, b => ci, o => s);
   and_1 : and2_312 port map( a => a, b => b, o => s2);
   and_2 : and2_311 port map( a => s1, b => ci, o => s3);
   or_1 : or2_154 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_153 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_153;

architecture SYN_Structural of fa_153 is

   component or2_153
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_309
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_310
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_309
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_310
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_310 port map( a => a, b => b, o => s1);
   xor_2 : xor2_309 port map( a => s1, b => ci, o => s);
   and_1 : and2_310 port map( a => a, b => b, o => s2);
   and_2 : and2_309 port map( a => s1, b => ci, o => s3);
   or_1 : or2_153 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_152 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_152;

architecture SYN_Structural of fa_152 is

   component or2_152
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_307
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_308
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_307
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_308
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_308 port map( a => a, b => b, o => s1);
   xor_2 : xor2_307 port map( a => s1, b => ci, o => s);
   and_1 : and2_308 port map( a => a, b => b, o => s2);
   and_2 : and2_307 port map( a => s1, b => ci, o => s3);
   or_1 : or2_152 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_151 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_151;

architecture SYN_Structural of fa_151 is

   component or2_151
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_305
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_306
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_305
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_306
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_306 port map( a => a, b => b, o => s1);
   xor_2 : xor2_305 port map( a => s1, b => ci, o => s);
   and_1 : and2_306 port map( a => a, b => b, o => s2);
   and_2 : and2_305 port map( a => s1, b => ci, o => s3);
   or_1 : or2_151 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_150 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_150;

architecture SYN_Structural of fa_150 is

   component or2_150
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_303
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_304
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_303
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_304
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_304 port map( a => a, b => b, o => s1);
   xor_2 : xor2_303 port map( a => s1, b => ci, o => s);
   and_1 : and2_304 port map( a => a, b => b, o => s2);
   and_2 : and2_303 port map( a => s1, b => ci, o => s3);
   or_1 : or2_150 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_149 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_149;

architecture SYN_Structural of fa_149 is

   component or2_149
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_301
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_302
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_301
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_302
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_302 port map( a => a, b => b, o => s1);
   xor_2 : xor2_301 port map( a => s1, b => ci, o => s);
   and_1 : and2_302 port map( a => a, b => b, o => s2);
   and_2 : and2_301 port map( a => s1, b => ci, o => s3);
   or_1 : or2_149 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_148 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_148;

architecture SYN_Structural of fa_148 is

   component or2_148
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_299
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_300
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_299
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_300
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_300 port map( a => a, b => b, o => s1);
   xor_2 : xor2_299 port map( a => s1, b => ci, o => s);
   and_1 : and2_300 port map( a => a, b => b, o => s2);
   and_2 : and2_299 port map( a => s1, b => ci, o => s3);
   or_1 : or2_148 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_147 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_147;

architecture SYN_Structural of fa_147 is

   component or2_147
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_297
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_298
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_297
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_298
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_298 port map( a => a, b => b, o => s1);
   xor_2 : xor2_297 port map( a => s1, b => ci, o => s);
   and_1 : and2_298 port map( a => a, b => b, o => s2);
   and_2 : and2_297 port map( a => s1, b => ci, o => s3);
   or_1 : or2_147 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_146 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_146;

architecture SYN_Structural of fa_146 is

   component or2_146
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_295
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_296
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_295
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_296
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_296 port map( a => a, b => b, o => s1);
   xor_2 : xor2_295 port map( a => s1, b => ci, o => s);
   and_1 : and2_296 port map( a => a, b => b, o => s2);
   and_2 : and2_295 port map( a => s1, b => ci, o => s3);
   or_1 : or2_146 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_145 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_145;

architecture SYN_Structural of fa_145 is

   component or2_145
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_293
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_294
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_293
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_294
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_294 port map( a => a, b => b, o => s1);
   xor_2 : xor2_293 port map( a => s1, b => ci, o => s);
   and_1 : and2_294 port map( a => a, b => b, o => s2);
   and_2 : and2_293 port map( a => s1, b => ci, o => s3);
   or_1 : or2_145 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_144 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_144;

architecture SYN_Structural of fa_144 is

   component or2_144
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_291
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_292
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_291
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_292
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_292 port map( a => a, b => b, o => s1);
   xor_2 : xor2_291 port map( a => s1, b => ci, o => s);
   and_1 : and2_292 port map( a => a, b => b, o => s2);
   and_2 : and2_291 port map( a => s1, b => ci, o => s3);
   or_1 : or2_144 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_143 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_143;

architecture SYN_Structural of fa_143 is

   component or2_143
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_289
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_290
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_289
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_290
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_290 port map( a => a, b => b, o => s1);
   xor_2 : xor2_289 port map( a => s1, b => ci, o => s);
   and_1 : and2_290 port map( a => a, b => b, o => s2);
   and_2 : and2_289 port map( a => s1, b => ci, o => s3);
   or_1 : or2_143 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_142 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_142;

architecture SYN_Structural of fa_142 is

   component or2_142
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_287
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_288
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_287
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_288
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_288 port map( a => a, b => b, o => s1);
   xor_2 : xor2_287 port map( a => s1, b => ci, o => s);
   and_1 : and2_288 port map( a => a, b => b, o => s2);
   and_2 : and2_287 port map( a => s1, b => ci, o => s3);
   or_1 : or2_142 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_141 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_141;

architecture SYN_Structural of fa_141 is

   component or2_141
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_285
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_286
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_285
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_286
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_286 port map( a => a, b => b, o => s1);
   xor_2 : xor2_285 port map( a => s1, b => ci, o => s);
   and_1 : and2_286 port map( a => a, b => b, o => s2);
   and_2 : and2_285 port map( a => s1, b => ci, o => s3);
   or_1 : or2_141 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_140 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_140;

architecture SYN_Structural of fa_140 is

   component or2_140
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_283
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_284
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_283
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_284
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_284 port map( a => a, b => b, o => s1);
   xor_2 : xor2_283 port map( a => s1, b => ci, o => s);
   and_1 : and2_284 port map( a => a, b => b, o => s2);
   and_2 : and2_283 port map( a => s1, b => ci, o => s3);
   or_1 : or2_140 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_139 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_139;

architecture SYN_Structural of fa_139 is

   component or2_139
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_281
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_282
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_281
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_282
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_282 port map( a => a, b => b, o => s1);
   xor_2 : xor2_281 port map( a => s1, b => ci, o => s);
   and_1 : and2_282 port map( a => a, b => b, o => s2);
   and_2 : and2_281 port map( a => s1, b => ci, o => s3);
   or_1 : or2_139 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_138 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_138;

architecture SYN_Structural of fa_138 is

   component or2_138
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_279
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_280
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_279
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_280
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_280 port map( a => a, b => b, o => s1);
   xor_2 : xor2_279 port map( a => s1, b => ci, o => s);
   and_1 : and2_280 port map( a => a, b => b, o => s2);
   and_2 : and2_279 port map( a => s1, b => ci, o => s3);
   or_1 : or2_138 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_137 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_137;

architecture SYN_Structural of fa_137 is

   component or2_137
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_277
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_278
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_277
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_278
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_278 port map( a => a, b => b, o => s1);
   xor_2 : xor2_277 port map( a => s1, b => ci, o => s);
   and_1 : and2_278 port map( a => a, b => b, o => s2);
   and_2 : and2_277 port map( a => s1, b => ci, o => s3);
   or_1 : or2_137 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_136 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_136;

architecture SYN_Structural of fa_136 is

   component or2_136
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_275
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_276
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_275
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_276
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_276 port map( a => a, b => b, o => s1);
   xor_2 : xor2_275 port map( a => s1, b => ci, o => s);
   and_1 : and2_276 port map( a => a, b => b, o => s2);
   and_2 : and2_275 port map( a => s1, b => ci, o => s3);
   or_1 : or2_136 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_135 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_135;

architecture SYN_Structural of fa_135 is

   component or2_135
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_273
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_274
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_273
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_274
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_274 port map( a => a, b => b, o => s1);
   xor_2 : xor2_273 port map( a => s1, b => ci, o => s);
   and_1 : and2_274 port map( a => a, b => b, o => s2);
   and_2 : and2_273 port map( a => s1, b => ci, o => s3);
   or_1 : or2_135 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_134 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_134;

architecture SYN_Structural of fa_134 is

   component or2_134
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_271
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_272
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_271
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_272
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_272 port map( a => a, b => b, o => s1);
   xor_2 : xor2_271 port map( a => s1, b => ci, o => s);
   and_1 : and2_272 port map( a => a, b => b, o => s2);
   and_2 : and2_271 port map( a => s1, b => ci, o => s3);
   or_1 : or2_134 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_133 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_133;

architecture SYN_Structural of fa_133 is

   component or2_133
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_269
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_270
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_269
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_270
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_270 port map( a => a, b => b, o => s1);
   xor_2 : xor2_269 port map( a => s1, b => ci, o => s);
   and_1 : and2_270 port map( a => a, b => b, o => s2);
   and_2 : and2_269 port map( a => s1, b => ci, o => s3);
   or_1 : or2_133 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_132 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_132;

architecture SYN_Structural of fa_132 is

   component or2_132
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_267
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_268
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_267
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_268
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_268 port map( a => a, b => b, o => s1);
   xor_2 : xor2_267 port map( a => s1, b => ci, o => s);
   and_1 : and2_268 port map( a => a, b => b, o => s2);
   and_2 : and2_267 port map( a => s1, b => ci, o => s3);
   or_1 : or2_132 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_131 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_131;

architecture SYN_Structural of fa_131 is

   component or2_131
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_265
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_266
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_265
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_266
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_266 port map( a => a, b => b, o => s1);
   xor_2 : xor2_265 port map( a => s1, b => ci, o => s);
   and_1 : and2_266 port map( a => a, b => b, o => s2);
   and_2 : and2_265 port map( a => s1, b => ci, o => s3);
   or_1 : or2_131 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_130 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_130;

architecture SYN_Structural of fa_130 is

   component or2_130
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_263
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_264
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_263
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_264
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_264 port map( a => a, b => b, o => s1);
   xor_2 : xor2_263 port map( a => s1, b => ci, o => s);
   and_1 : and2_264 port map( a => a, b => b, o => s2);
   and_2 : and2_263 port map( a => s1, b => ci, o => s3);
   or_1 : or2_130 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_129 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_129;

architecture SYN_Structural of fa_129 is

   component or2_129
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_261
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_262
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_261
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_262
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_262 port map( a => a, b => b, o => s1);
   xor_2 : xor2_261 port map( a => s1, b => ci, o => s);
   and_1 : and2_262 port map( a => a, b => b, o => s2);
   and_2 : and2_261 port map( a => s1, b => ci, o => s3);
   or_1 : or2_129 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_128 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_128;

architecture SYN_Structural of fa_128 is

   component or2_128
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_259
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_260
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_259
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_260
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_260 port map( a => a, b => b, o => s1);
   xor_2 : xor2_259 port map( a => s1, b => ci, o => s);
   and_1 : and2_260 port map( a => a, b => b, o => s2);
   and_2 : and2_259 port map( a => s1, b => ci, o => s3);
   or_1 : or2_128 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_127 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_127;

architecture SYN_Structural of fa_127 is

   component or2_127
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_257
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_258
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_257
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_258
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_258 port map( a => a, b => b, o => s1);
   xor_2 : xor2_257 port map( a => s1, b => ci, o => s);
   and_1 : and2_258 port map( a => a, b => b, o => s2);
   and_2 : and2_257 port map( a => s1, b => ci, o => s3);
   or_1 : or2_127 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_126 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_126;

architecture SYN_Structural of fa_126 is

   component or2_126
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_255
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_256
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_255
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_256
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_256 port map( a => a, b => b, o => s1);
   xor_2 : xor2_255 port map( a => s1, b => ci, o => s);
   and_1 : and2_256 port map( a => a, b => b, o => s2);
   and_2 : and2_255 port map( a => s1, b => ci, o => s3);
   or_1 : or2_126 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_125 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_125;

architecture SYN_Structural of fa_125 is

   component or2_125
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_253
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_254
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_253
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_254
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_254 port map( a => a, b => b, o => s1);
   xor_2 : xor2_253 port map( a => s1, b => ci, o => s);
   and_1 : and2_254 port map( a => a, b => b, o => s2);
   and_2 : and2_253 port map( a => s1, b => ci, o => s3);
   or_1 : or2_125 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_124 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_124;

architecture SYN_Structural of fa_124 is

   component or2_124
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_250
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_251
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_250
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_251
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_251 port map( a => a, b => b, o => s1);
   xor_2 : xor2_250 port map( a => s1, b => ci, o => s);
   and_1 : and2_251 port map( a => a, b => b, o => s2);
   and_2 : and2_250 port map( a => s1, b => ci, o => s3);
   or_1 : or2_124 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_123 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_123;

architecture SYN_Structural of fa_123 is

   component or2_123
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_248
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_249
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_248
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_249
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_249 port map( a => a, b => b, o => s1);
   xor_2 : xor2_248 port map( a => s1, b => ci, o => s);
   and_1 : and2_249 port map( a => a, b => b, o => s2);
   and_2 : and2_248 port map( a => s1, b => ci, o => s3);
   or_1 : or2_123 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_122 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_122;

architecture SYN_Structural of fa_122 is

   component or2_122
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_246
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_247
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_246
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_247
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_247 port map( a => a, b => b, o => s1);
   xor_2 : xor2_246 port map( a => s1, b => ci, o => s);
   and_1 : and2_247 port map( a => a, b => b, o => s2);
   and_2 : and2_246 port map( a => s1, b => ci, o => s3);
   or_1 : or2_122 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_121 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_121;

architecture SYN_Structural of fa_121 is

   component or2_121
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_244
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_245
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_244
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_245
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_245 port map( a => a, b => b, o => s1);
   xor_2 : xor2_244 port map( a => s1, b => ci, o => s);
   and_1 : and2_245 port map( a => a, b => b, o => s2);
   and_2 : and2_244 port map( a => s1, b => ci, o => s3);
   or_1 : or2_121 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_120 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_120;

architecture SYN_Structural of fa_120 is

   component or2_120
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_242
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_243
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_242
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_243
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_243 port map( a => a, b => b, o => s1);
   xor_2 : xor2_242 port map( a => s1, b => ci, o => s);
   and_1 : and2_243 port map( a => a, b => b, o => s2);
   and_2 : and2_242 port map( a => s1, b => ci, o => s3);
   or_1 : or2_120 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_119 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_119;

architecture SYN_Structural of fa_119 is

   component or2_119
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_240
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_241
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_240
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_241
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_241 port map( a => a, b => b, o => s1);
   xor_2 : xor2_240 port map( a => s1, b => ci, o => s);
   and_1 : and2_241 port map( a => a, b => b, o => s2);
   and_2 : and2_240 port map( a => s1, b => ci, o => s3);
   or_1 : or2_119 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_118 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_118;

architecture SYN_Structural of fa_118 is

   component or2_118
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_238
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_239
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_238
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_239
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_239 port map( a => a, b => b, o => s1);
   xor_2 : xor2_238 port map( a => s1, b => ci, o => s);
   and_1 : and2_239 port map( a => a, b => b, o => s2);
   and_2 : and2_238 port map( a => s1, b => ci, o => s3);
   or_1 : or2_118 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_117 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_117;

architecture SYN_Structural of fa_117 is

   component or2_117
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_236
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_237
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_236
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_237
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_237 port map( a => a, b => b, o => s1);
   xor_2 : xor2_236 port map( a => s1, b => ci, o => s);
   and_1 : and2_237 port map( a => a, b => b, o => s2);
   and_2 : and2_236 port map( a => s1, b => ci, o => s3);
   or_1 : or2_117 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_116 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_116;

architecture SYN_Structural of fa_116 is

   component or2_116
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_234
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_235
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_234
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_235
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_235 port map( a => a, b => b, o => s1);
   xor_2 : xor2_234 port map( a => s1, b => ci, o => s);
   and_1 : and2_235 port map( a => a, b => b, o => s2);
   and_2 : and2_234 port map( a => s1, b => ci, o => s3);
   or_1 : or2_116 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_115 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_115;

architecture SYN_Structural of fa_115 is

   component or2_115
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_232
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_233
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_232
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_233
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_233 port map( a => a, b => b, o => s1);
   xor_2 : xor2_232 port map( a => s1, b => ci, o => s);
   and_1 : and2_233 port map( a => a, b => b, o => s2);
   and_2 : and2_232 port map( a => s1, b => ci, o => s3);
   or_1 : or2_115 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_114 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_114;

architecture SYN_Structural of fa_114 is

   component or2_114
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_230
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_231
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_230
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_231
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_231 port map( a => a, b => b, o => s1);
   xor_2 : xor2_230 port map( a => s1, b => ci, o => s);
   and_1 : and2_231 port map( a => a, b => b, o => s2);
   and_2 : and2_230 port map( a => s1, b => ci, o => s3);
   or_1 : or2_114 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_113 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_113;

architecture SYN_Structural of fa_113 is

   component or2_113
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_228
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_229
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_228
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_229
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_229 port map( a => a, b => b, o => s1);
   xor_2 : xor2_228 port map( a => s1, b => ci, o => s);
   and_1 : and2_229 port map( a => a, b => b, o => s2);
   and_2 : and2_228 port map( a => s1, b => ci, o => s3);
   or_1 : or2_113 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_112 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_112;

architecture SYN_Structural of fa_112 is

   component or2_112
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_226
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_227
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_226
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_227
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_227 port map( a => a, b => b, o => s1);
   xor_2 : xor2_226 port map( a => s1, b => ci, o => s);
   and_1 : and2_227 port map( a => a, b => b, o => s2);
   and_2 : and2_226 port map( a => s1, b => ci, o => s3);
   or_1 : or2_112 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_111 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_111;

architecture SYN_Structural of fa_111 is

   component or2_111
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_224
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_225
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_224
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_225
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_225 port map( a => a, b => b, o => s1);
   xor_2 : xor2_224 port map( a => s1, b => ci, o => s);
   and_1 : and2_225 port map( a => a, b => b, o => s2);
   and_2 : and2_224 port map( a => s1, b => ci, o => s3);
   or_1 : or2_111 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_110 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_110;

architecture SYN_Structural of fa_110 is

   component or2_110
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_222
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_223
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_222
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_223
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_223 port map( a => a, b => b, o => s1);
   xor_2 : xor2_222 port map( a => s1, b => ci, o => s);
   and_1 : and2_223 port map( a => a, b => b, o => s2);
   and_2 : and2_222 port map( a => s1, b => ci, o => s3);
   or_1 : or2_110 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_109 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_109;

architecture SYN_Structural of fa_109 is

   component or2_109
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_220
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_221
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_220
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_221
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_221 port map( a => a, b => b, o => s1);
   xor_2 : xor2_220 port map( a => s1, b => ci, o => s);
   and_1 : and2_221 port map( a => a, b => b, o => s2);
   and_2 : and2_220 port map( a => s1, b => ci, o => s3);
   or_1 : or2_109 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_108 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_108;

architecture SYN_Structural of fa_108 is

   component or2_108
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_218
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_219
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_218
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_219
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_219 port map( a => a, b => b, o => s1);
   xor_2 : xor2_218 port map( a => s1, b => ci, o => s);
   and_1 : and2_219 port map( a => a, b => b, o => s2);
   and_2 : and2_218 port map( a => s1, b => ci, o => s3);
   or_1 : or2_108 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_107 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_107;

architecture SYN_Structural of fa_107 is

   component or2_107
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_216
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_217
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_216
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_217
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_217 port map( a => a, b => b, o => s1);
   xor_2 : xor2_216 port map( a => s1, b => ci, o => s);
   and_1 : and2_217 port map( a => a, b => b, o => s2);
   and_2 : and2_216 port map( a => s1, b => ci, o => s3);
   or_1 : or2_107 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_106 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_106;

architecture SYN_Structural of fa_106 is

   component or2_106
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_214
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_215
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_214
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_215
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_215 port map( a => a, b => b, o => s1);
   xor_2 : xor2_214 port map( a => s1, b => ci, o => s);
   and_1 : and2_215 port map( a => a, b => b, o => s2);
   and_2 : and2_214 port map( a => s1, b => ci, o => s3);
   or_1 : or2_106 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_105 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_105;

architecture SYN_Structural of fa_105 is

   component or2_105
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_212
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_213
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_212
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_213
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_213 port map( a => a, b => b, o => s1);
   xor_2 : xor2_212 port map( a => s1, b => ci, o => s);
   and_1 : and2_213 port map( a => a, b => b, o => s2);
   and_2 : and2_212 port map( a => s1, b => ci, o => s3);
   or_1 : or2_105 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_104 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_104;

architecture SYN_Structural of fa_104 is

   component or2_104
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_210
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_211
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_210
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_211
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_211 port map( a => a, b => b, o => s1);
   xor_2 : xor2_210 port map( a => s1, b => ci, o => s);
   and_1 : and2_211 port map( a => a, b => b, o => s2);
   and_2 : and2_210 port map( a => s1, b => ci, o => s3);
   or_1 : or2_104 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_103 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_103;

architecture SYN_Structural of fa_103 is

   component or2_103
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_208
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_209
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_208
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_209
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_209 port map( a => a, b => b, o => s1);
   xor_2 : xor2_208 port map( a => s1, b => ci, o => s);
   and_1 : and2_209 port map( a => a, b => b, o => s2);
   and_2 : and2_208 port map( a => s1, b => ci, o => s3);
   or_1 : or2_103 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_102 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_102;

architecture SYN_Structural of fa_102 is

   component or2_102
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_206
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_207
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_206
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_207
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_207 port map( a => a, b => b, o => s1);
   xor_2 : xor2_206 port map( a => s1, b => ci, o => s);
   and_1 : and2_207 port map( a => a, b => b, o => s2);
   and_2 : and2_206 port map( a => s1, b => ci, o => s3);
   or_1 : or2_102 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_101 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_101;

architecture SYN_Structural of fa_101 is

   component or2_101
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_204
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_205
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_204
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_205
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_205 port map( a => a, b => b, o => s1);
   xor_2 : xor2_204 port map( a => s1, b => ci, o => s);
   and_1 : and2_205 port map( a => a, b => b, o => s2);
   and_2 : and2_204 port map( a => s1, b => ci, o => s3);
   or_1 : or2_101 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_100 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_100;

architecture SYN_Structural of fa_100 is

   component or2_100
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_202
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_203
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_202
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_203
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_203 port map( a => a, b => b, o => s1);
   xor_2 : xor2_202 port map( a => s1, b => ci, o => s);
   and_1 : and2_203 port map( a => a, b => b, o => s2);
   and_2 : and2_202 port map( a => s1, b => ci, o => s3);
   or_1 : or2_100 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_99 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_99;

architecture SYN_Structural of fa_99 is

   component or2_99
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_200
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_201
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_200
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_201
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_201 port map( a => a, b => b, o => s1);
   xor_2 : xor2_200 port map( a => s1, b => ci, o => s);
   and_1 : and2_201 port map( a => a, b => b, o => s2);
   and_2 : and2_200 port map( a => s1, b => ci, o => s3);
   or_1 : or2_99 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_98 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_98;

architecture SYN_Structural of fa_98 is

   component or2_98
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_198
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_199
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_198
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_199
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_199 port map( a => a, b => b, o => s1);
   xor_2 : xor2_198 port map( a => s1, b => ci, o => s);
   and_1 : and2_199 port map( a => a, b => b, o => s2);
   and_2 : and2_198 port map( a => s1, b => ci, o => s3);
   or_1 : or2_98 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_97 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_97;

architecture SYN_Structural of fa_97 is

   component or2_97
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_196
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_197
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_196
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_197
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_197 port map( a => a, b => b, o => s1);
   xor_2 : xor2_196 port map( a => s1, b => ci, o => s);
   and_1 : and2_197 port map( a => a, b => b, o => s2);
   and_2 : and2_196 port map( a => s1, b => ci, o => s3);
   or_1 : or2_97 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_96 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_96;

architecture SYN_Structural of fa_96 is

   component or2_96
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_194
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_195
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_194
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_195
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_195 port map( a => a, b => b, o => s1);
   xor_2 : xor2_194 port map( a => s1, b => ci, o => s);
   and_1 : and2_195 port map( a => a, b => b, o => s2);
   and_2 : and2_194 port map( a => s1, b => ci, o => s3);
   or_1 : or2_96 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_95 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_95;

architecture SYN_Structural of fa_95 is

   component or2_95
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_192
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_193
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_192
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_193
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_193 port map( a => a, b => b, o => s1);
   xor_2 : xor2_192 port map( a => s1, b => ci, o => s);
   and_1 : and2_193 port map( a => a, b => b, o => s2);
   and_2 : and2_192 port map( a => s1, b => ci, o => s3);
   or_1 : or2_95 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_94 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_94;

architecture SYN_Structural of fa_94 is

   component or2_94
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_190
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_191
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_190
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_191
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_191 port map( a => a, b => b, o => s1);
   xor_2 : xor2_190 port map( a => s1, b => ci, o => s);
   and_1 : and2_191 port map( a => a, b => b, o => s2);
   and_2 : and2_190 port map( a => s1, b => ci, o => s3);
   or_1 : or2_94 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_93 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_93;

architecture SYN_Structural of fa_93 is

   component or2_93
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_187
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_188
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_187
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_188
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_188 port map( a => a, b => b, o => s1);
   xor_2 : xor2_187 port map( a => s1, b => ci, o => s);
   and_1 : and2_188 port map( a => a, b => b, o => s2);
   and_2 : and2_187 port map( a => s1, b => ci, o => s3);
   or_1 : or2_93 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_92 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_92;

architecture SYN_Structural of fa_92 is

   component or2_92
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_185
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_186
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_185
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_186
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_186 port map( a => a, b => b, o => s1);
   xor_2 : xor2_185 port map( a => s1, b => ci, o => s);
   and_1 : and2_186 port map( a => a, b => b, o => s2);
   and_2 : and2_185 port map( a => s1, b => ci, o => s3);
   or_1 : or2_92 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_91 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_91;

architecture SYN_Structural of fa_91 is

   component or2_91
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_183
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_184
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_183
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_184
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_184 port map( a => a, b => b, o => s1);
   xor_2 : xor2_183 port map( a => s1, b => ci, o => s);
   and_1 : and2_184 port map( a => a, b => b, o => s2);
   and_2 : and2_183 port map( a => s1, b => ci, o => s3);
   or_1 : or2_91 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_90 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_90;

architecture SYN_Structural of fa_90 is

   component or2_90
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_181
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_182
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_181
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_182
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_182 port map( a => a, b => b, o => s1);
   xor_2 : xor2_181 port map( a => s1, b => ci, o => s);
   and_1 : and2_182 port map( a => a, b => b, o => s2);
   and_2 : and2_181 port map( a => s1, b => ci, o => s3);
   or_1 : or2_90 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_89 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_89;

architecture SYN_Structural of fa_89 is

   component or2_89
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_179
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_180
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_179
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_180
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_180 port map( a => a, b => b, o => s1);
   xor_2 : xor2_179 port map( a => s1, b => ci, o => s);
   and_1 : and2_180 port map( a => a, b => b, o => s2);
   and_2 : and2_179 port map( a => s1, b => ci, o => s3);
   or_1 : or2_89 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_88 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_88;

architecture SYN_Structural of fa_88 is

   component or2_88
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_177
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_178
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_177
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_178
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_178 port map( a => a, b => b, o => s1);
   xor_2 : xor2_177 port map( a => s1, b => ci, o => s);
   and_1 : and2_178 port map( a => a, b => b, o => s2);
   and_2 : and2_177 port map( a => s1, b => ci, o => s3);
   or_1 : or2_88 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_87 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_87;

architecture SYN_Structural of fa_87 is

   component or2_87
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_175
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_176
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_175
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_176
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_176 port map( a => a, b => b, o => s1);
   xor_2 : xor2_175 port map( a => s1, b => ci, o => s);
   and_1 : and2_176 port map( a => a, b => b, o => s2);
   and_2 : and2_175 port map( a => s1, b => ci, o => s3);
   or_1 : or2_87 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_86 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_86;

architecture SYN_Structural of fa_86 is

   component or2_86
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_173
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_174
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_173
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_174
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_174 port map( a => a, b => b, o => s1);
   xor_2 : xor2_173 port map( a => s1, b => ci, o => s);
   and_1 : and2_174 port map( a => a, b => b, o => s2);
   and_2 : and2_173 port map( a => s1, b => ci, o => s3);
   or_1 : or2_86 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_85 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_85;

architecture SYN_Structural of fa_85 is

   component or2_85
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_171
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_172
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_171
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_172
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_172 port map( a => a, b => b, o => s1);
   xor_2 : xor2_171 port map( a => s1, b => ci, o => s);
   and_1 : and2_172 port map( a => a, b => b, o => s2);
   and_2 : and2_171 port map( a => s1, b => ci, o => s3);
   or_1 : or2_85 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_84 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_84;

architecture SYN_Structural of fa_84 is

   component or2_84
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_169
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_170
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_169
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_170
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_170 port map( a => a, b => b, o => s1);
   xor_2 : xor2_169 port map( a => s1, b => ci, o => s);
   and_1 : and2_170 port map( a => a, b => b, o => s2);
   and_2 : and2_169 port map( a => s1, b => ci, o => s3);
   or_1 : or2_84 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_83 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_83;

architecture SYN_Structural of fa_83 is

   component or2_83
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_167
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_168
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_167
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_168
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_168 port map( a => a, b => b, o => s1);
   xor_2 : xor2_167 port map( a => s1, b => ci, o => s);
   and_1 : and2_168 port map( a => a, b => b, o => s2);
   and_2 : and2_167 port map( a => s1, b => ci, o => s3);
   or_1 : or2_83 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_82 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_82;

architecture SYN_Structural of fa_82 is

   component or2_82
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_165
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_166
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_165
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_166
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_166 port map( a => a, b => b, o => s1);
   xor_2 : xor2_165 port map( a => s1, b => ci, o => s);
   and_1 : and2_166 port map( a => a, b => b, o => s2);
   and_2 : and2_165 port map( a => s1, b => ci, o => s3);
   or_1 : or2_82 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_81 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_81;

architecture SYN_Structural of fa_81 is

   component or2_81
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_163
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_164
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_163
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_164
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_164 port map( a => a, b => b, o => s1);
   xor_2 : xor2_163 port map( a => s1, b => ci, o => s);
   and_1 : and2_164 port map( a => a, b => b, o => s2);
   and_2 : and2_163 port map( a => s1, b => ci, o => s3);
   or_1 : or2_81 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_80 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_80;

architecture SYN_Structural of fa_80 is

   component or2_80
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_161
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_162
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_161
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_162
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_162 port map( a => a, b => b, o => s1);
   xor_2 : xor2_161 port map( a => s1, b => ci, o => s);
   and_1 : and2_162 port map( a => a, b => b, o => s2);
   and_2 : and2_161 port map( a => s1, b => ci, o => s3);
   or_1 : or2_80 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_79 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_79;

architecture SYN_Structural of fa_79 is

   component or2_79
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_159
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_160
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_159
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_160
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_160 port map( a => a, b => b, o => s1);
   xor_2 : xor2_159 port map( a => s1, b => ci, o => s);
   and_1 : and2_160 port map( a => a, b => b, o => s2);
   and_2 : and2_159 port map( a => s1, b => ci, o => s3);
   or_1 : or2_79 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_78 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_78;

architecture SYN_Structural of fa_78 is

   component or2_78
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_157
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_158
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_157
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_158
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_158 port map( a => a, b => b, o => s1);
   xor_2 : xor2_157 port map( a => s1, b => ci, o => s);
   and_1 : and2_158 port map( a => a, b => b, o => s2);
   and_2 : and2_157 port map( a => s1, b => ci, o => s3);
   or_1 : or2_78 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_77 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_77;

architecture SYN_Structural of fa_77 is

   component or2_77
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_155
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_156
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_155
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_156
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_156 port map( a => a, b => b, o => s1);
   xor_2 : xor2_155 port map( a => s1, b => ci, o => s);
   and_1 : and2_156 port map( a => a, b => b, o => s2);
   and_2 : and2_155 port map( a => s1, b => ci, o => s3);
   or_1 : or2_77 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_76 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_76;

architecture SYN_Structural of fa_76 is

   component or2_76
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_153
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_154
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_153
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_154
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_154 port map( a => a, b => b, o => s1);
   xor_2 : xor2_153 port map( a => s1, b => ci, o => s);
   and_1 : and2_154 port map( a => a, b => b, o => s2);
   and_2 : and2_153 port map( a => s1, b => ci, o => s3);
   or_1 : or2_76 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_75 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_75;

architecture SYN_Structural of fa_75 is

   component or2_75
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_151
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_152
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_151
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_152
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_152 port map( a => a, b => b, o => s1);
   xor_2 : xor2_151 port map( a => s1, b => ci, o => s);
   and_1 : and2_152 port map( a => a, b => b, o => s2);
   and_2 : and2_151 port map( a => s1, b => ci, o => s3);
   or_1 : or2_75 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_74 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_74;

architecture SYN_Structural of fa_74 is

   component or2_74
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_149
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_150
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_149
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_150
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_150 port map( a => a, b => b, o => s1);
   xor_2 : xor2_149 port map( a => s1, b => ci, o => s);
   and_1 : and2_150 port map( a => a, b => b, o => s2);
   and_2 : and2_149 port map( a => s1, b => ci, o => s3);
   or_1 : or2_74 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_73 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_73;

architecture SYN_Structural of fa_73 is

   component or2_73
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_147
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_148
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_147
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_148
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_148 port map( a => a, b => b, o => s1);
   xor_2 : xor2_147 port map( a => s1, b => ci, o => s);
   and_1 : and2_148 port map( a => a, b => b, o => s2);
   and_2 : and2_147 port map( a => s1, b => ci, o => s3);
   or_1 : or2_73 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_72 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_72;

architecture SYN_Structural of fa_72 is

   component or2_72
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_145
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_146
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_145
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_146
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_146 port map( a => a, b => b, o => s1);
   xor_2 : xor2_145 port map( a => s1, b => ci, o => s);
   and_1 : and2_146 port map( a => a, b => b, o => s2);
   and_2 : and2_145 port map( a => s1, b => ci, o => s3);
   or_1 : or2_72 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_71 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_71;

architecture SYN_Structural of fa_71 is

   component or2_71
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_143
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_144
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_143
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_144
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_144 port map( a => a, b => b, o => s1);
   xor_2 : xor2_143 port map( a => s1, b => ci, o => s);
   and_1 : and2_144 port map( a => a, b => b, o => s2);
   and_2 : and2_143 port map( a => s1, b => ci, o => s3);
   or_1 : or2_71 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_70 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_70;

architecture SYN_Structural of fa_70 is

   component or2_70
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_141
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_142
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_141
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_142
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_142 port map( a => a, b => b, o => s1);
   xor_2 : xor2_141 port map( a => s1, b => ci, o => s);
   and_1 : and2_142 port map( a => a, b => b, o => s2);
   and_2 : and2_141 port map( a => s1, b => ci, o => s3);
   or_1 : or2_70 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_69 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_69;

architecture SYN_Structural of fa_69 is

   component or2_69
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_139
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_140
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_139
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_140
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_140 port map( a => a, b => b, o => s1);
   xor_2 : xor2_139 port map( a => s1, b => ci, o => s);
   and_1 : and2_140 port map( a => a, b => b, o => s2);
   and_2 : and2_139 port map( a => s1, b => ci, o => s3);
   or_1 : or2_69 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_68 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_68;

architecture SYN_Structural of fa_68 is

   component or2_68
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_137
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_138
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_137
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_138
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_138 port map( a => a, b => b, o => s1);
   xor_2 : xor2_137 port map( a => s1, b => ci, o => s);
   and_1 : and2_138 port map( a => a, b => b, o => s2);
   and_2 : and2_137 port map( a => s1, b => ci, o => s3);
   or_1 : or2_68 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_67 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_67;

architecture SYN_Structural of fa_67 is

   component or2_67
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_135
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_136
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_135
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_136
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_136 port map( a => a, b => b, o => s1);
   xor_2 : xor2_135 port map( a => s1, b => ci, o => s);
   and_1 : and2_136 port map( a => a, b => b, o => s2);
   and_2 : and2_135 port map( a => s1, b => ci, o => s3);
   or_1 : or2_67 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_66 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_66;

architecture SYN_Structural of fa_66 is

   component or2_66
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_133
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_134
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_133
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_134
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_134 port map( a => a, b => b, o => s1);
   xor_2 : xor2_133 port map( a => s1, b => ci, o => s);
   and_1 : and2_134 port map( a => a, b => b, o => s2);
   and_2 : and2_133 port map( a => s1, b => ci, o => s3);
   or_1 : or2_66 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_65 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_65;

architecture SYN_Structural of fa_65 is

   component or2_65
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_131
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_132
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_131
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_132
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_132 port map( a => a, b => b, o => s1);
   xor_2 : xor2_131 port map( a => s1, b => ci, o => s);
   and_1 : and2_132 port map( a => a, b => b, o => s2);
   and_2 : and2_131 port map( a => s1, b => ci, o => s3);
   or_1 : or2_65 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_64 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_64;

architecture SYN_Structural of fa_64 is

   component or2_64
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_129
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_130
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_129
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_130
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_130 port map( a => a, b => b, o => s1);
   xor_2 : xor2_129 port map( a => s1, b => ci, o => s);
   and_1 : and2_130 port map( a => a, b => b, o => s2);
   and_2 : and2_129 port map( a => s1, b => ci, o => s3);
   or_1 : or2_64 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_63 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_63;

architecture SYN_Structural of fa_63 is

   component or2_63
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_127
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_128
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_127
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_128
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_128 port map( a => a, b => b, o => s1);
   xor_2 : xor2_127 port map( a => s1, b => ci, o => s);
   and_1 : and2_128 port map( a => a, b => b, o => s2);
   and_2 : and2_127 port map( a => s1, b => ci, o => s3);
   or_1 : or2_63 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_62 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_62;

architecture SYN_Structural of fa_62 is

   component or2_62
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_124
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_125
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_124
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_125
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_125 port map( a => a, b => b, o => s1);
   xor_2 : xor2_124 port map( a => s1, b => ci, o => s);
   and_1 : and2_125 port map( a => a, b => b, o => s2);
   and_2 : and2_124 port map( a => s1, b => ci, o => s3);
   or_1 : or2_62 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_61 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_61;

architecture SYN_Structural of fa_61 is

   component or2_61
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_122
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_123
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_122
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_123
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_123 port map( a => a, b => b, o => s1);
   xor_2 : xor2_122 port map( a => s1, b => ci, o => s);
   and_1 : and2_123 port map( a => a, b => b, o => s2);
   and_2 : and2_122 port map( a => s1, b => ci, o => s3);
   or_1 : or2_61 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_60 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_60;

architecture SYN_Structural of fa_60 is

   component or2_60
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_120
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_121
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_120
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_121
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_121 port map( a => a, b => b, o => s1);
   xor_2 : xor2_120 port map( a => s1, b => ci, o => s);
   and_1 : and2_121 port map( a => a, b => b, o => s2);
   and_2 : and2_120 port map( a => s1, b => ci, o => s3);
   or_1 : or2_60 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_59 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_59;

architecture SYN_Structural of fa_59 is

   component or2_59
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_118
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_119
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_118
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_119
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_119 port map( a => a, b => b, o => s1);
   xor_2 : xor2_118 port map( a => s1, b => ci, o => s);
   and_1 : and2_119 port map( a => a, b => b, o => s2);
   and_2 : and2_118 port map( a => s1, b => ci, o => s3);
   or_1 : or2_59 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_58 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_58;

architecture SYN_Structural of fa_58 is

   component or2_58
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_116
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_117
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_116
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_117
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_117 port map( a => a, b => b, o => s1);
   xor_2 : xor2_116 port map( a => s1, b => ci, o => s);
   and_1 : and2_117 port map( a => a, b => b, o => s2);
   and_2 : and2_116 port map( a => s1, b => ci, o => s3);
   or_1 : or2_58 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_57 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_57;

architecture SYN_Structural of fa_57 is

   component or2_57
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_114
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_115
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_114
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_115
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_115 port map( a => a, b => b, o => s1);
   xor_2 : xor2_114 port map( a => s1, b => ci, o => s);
   and_1 : and2_115 port map( a => a, b => b, o => s2);
   and_2 : and2_114 port map( a => s1, b => ci, o => s3);
   or_1 : or2_57 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_56 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_56;

architecture SYN_Structural of fa_56 is

   component or2_56
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_112
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_113
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_112
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_113
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_113 port map( a => a, b => b, o => s1);
   xor_2 : xor2_112 port map( a => s1, b => ci, o => s);
   and_1 : and2_113 port map( a => a, b => b, o => s2);
   and_2 : and2_112 port map( a => s1, b => ci, o => s3);
   or_1 : or2_56 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_55 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_55;

architecture SYN_Structural of fa_55 is

   component or2_55
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_110
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_111
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_110
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_111
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_111 port map( a => a, b => b, o => s1);
   xor_2 : xor2_110 port map( a => s1, b => ci, o => s);
   and_1 : and2_111 port map( a => a, b => b, o => s2);
   and_2 : and2_110 port map( a => s1, b => ci, o => s3);
   or_1 : or2_55 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_54 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_54;

architecture SYN_Structural of fa_54 is

   component or2_54
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_108
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_109
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_108
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_109
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_109 port map( a => a, b => b, o => s1);
   xor_2 : xor2_108 port map( a => s1, b => ci, o => s);
   and_1 : and2_109 port map( a => a, b => b, o => s2);
   and_2 : and2_108 port map( a => s1, b => ci, o => s3);
   or_1 : or2_54 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_53 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_53;

architecture SYN_Structural of fa_53 is

   component or2_53
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_106
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_107
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_106
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_107
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_107 port map( a => a, b => b, o => s1);
   xor_2 : xor2_106 port map( a => s1, b => ci, o => s);
   and_1 : and2_107 port map( a => a, b => b, o => s2);
   and_2 : and2_106 port map( a => s1, b => ci, o => s3);
   or_1 : or2_53 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_52 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_52;

architecture SYN_Structural of fa_52 is

   component or2_52
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_104
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_105
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_104
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_105
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_105 port map( a => a, b => b, o => s1);
   xor_2 : xor2_104 port map( a => s1, b => ci, o => s);
   and_1 : and2_105 port map( a => a, b => b, o => s2);
   and_2 : and2_104 port map( a => s1, b => ci, o => s3);
   or_1 : or2_52 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_51 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_51;

architecture SYN_Structural of fa_51 is

   component or2_51
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_102
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_103
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_102
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_103
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_103 port map( a => a, b => b, o => s1);
   xor_2 : xor2_102 port map( a => s1, b => ci, o => s);
   and_1 : and2_103 port map( a => a, b => b, o => s2);
   and_2 : and2_102 port map( a => s1, b => ci, o => s3);
   or_1 : or2_51 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_50 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_50;

architecture SYN_Structural of fa_50 is

   component or2_50
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_100
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_101
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_100
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_101
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_101 port map( a => a, b => b, o => s1);
   xor_2 : xor2_100 port map( a => s1, b => ci, o => s);
   and_1 : and2_101 port map( a => a, b => b, o => s2);
   and_2 : and2_100 port map( a => s1, b => ci, o => s3);
   or_1 : or2_50 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_49 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_49;

architecture SYN_Structural of fa_49 is

   component or2_49
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_98
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_99
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_98
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_99
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_99 port map( a => a, b => b, o => s1);
   xor_2 : xor2_98 port map( a => s1, b => ci, o => s);
   and_1 : and2_99 port map( a => a, b => b, o => s2);
   and_2 : and2_98 port map( a => s1, b => ci, o => s3);
   or_1 : or2_49 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_48 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_48;

architecture SYN_Structural of fa_48 is

   component or2_48
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_96
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_97
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_96
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_97
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_97 port map( a => a, b => b, o => s1);
   xor_2 : xor2_96 port map( a => s1, b => ci, o => s);
   and_1 : and2_97 port map( a => a, b => b, o => s2);
   and_2 : and2_96 port map( a => s1, b => ci, o => s3);
   or_1 : or2_48 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_47 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_47;

architecture SYN_Structural of fa_47 is

   component or2_47
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_94
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_95
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_94
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_95
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_95 port map( a => a, b => b, o => s1);
   xor_2 : xor2_94 port map( a => s1, b => ci, o => s);
   and_1 : and2_95 port map( a => a, b => b, o => s2);
   and_2 : and2_94 port map( a => s1, b => ci, o => s3);
   or_1 : or2_47 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_46 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_46;

architecture SYN_Structural of fa_46 is

   component or2_46
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_92
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_93
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_92
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_93
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_93 port map( a => a, b => b, o => s1);
   xor_2 : xor2_92 port map( a => s1, b => ci, o => s);
   and_1 : and2_93 port map( a => a, b => b, o => s2);
   and_2 : and2_92 port map( a => s1, b => ci, o => s3);
   or_1 : or2_46 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_45 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_45;

architecture SYN_Structural of fa_45 is

   component or2_45
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_90
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_91
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_90
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_91
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_91 port map( a => a, b => b, o => s1);
   xor_2 : xor2_90 port map( a => s1, b => ci, o => s);
   and_1 : and2_91 port map( a => a, b => b, o => s2);
   and_2 : and2_90 port map( a => s1, b => ci, o => s3);
   or_1 : or2_45 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_44 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_44;

architecture SYN_Structural of fa_44 is

   component or2_44
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_88
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_89
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_88
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_89
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_89 port map( a => a, b => b, o => s1);
   xor_2 : xor2_88 port map( a => s1, b => ci, o => s);
   and_1 : and2_89 port map( a => a, b => b, o => s2);
   and_2 : and2_88 port map( a => s1, b => ci, o => s3);
   or_1 : or2_44 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_43 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_43;

architecture SYN_Structural of fa_43 is

   component or2_43
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_86
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_87
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_86
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_87
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_87 port map( a => a, b => b, o => s1);
   xor_2 : xor2_86 port map( a => s1, b => ci, o => s);
   and_1 : and2_87 port map( a => a, b => b, o => s2);
   and_2 : and2_86 port map( a => s1, b => ci, o => s3);
   or_1 : or2_43 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_42 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_42;

architecture SYN_Structural of fa_42 is

   component or2_42
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_84
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_85
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_84
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_85
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_85 port map( a => a, b => b, o => s1);
   xor_2 : xor2_84 port map( a => s1, b => ci, o => s);
   and_1 : and2_85 port map( a => a, b => b, o => s2);
   and_2 : and2_84 port map( a => s1, b => ci, o => s3);
   or_1 : or2_42 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_41 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_41;

architecture SYN_Structural of fa_41 is

   component or2_41
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_82
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_83
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_82
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_83
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_83 port map( a => a, b => b, o => s1);
   xor_2 : xor2_82 port map( a => s1, b => ci, o => s);
   and_1 : and2_83 port map( a => a, b => b, o => s2);
   and_2 : and2_82 port map( a => s1, b => ci, o => s3);
   or_1 : or2_41 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_40 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_40;

architecture SYN_Structural of fa_40 is

   component or2_40
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_80
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_81
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_80
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_81
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_81 port map( a => a, b => b, o => s1);
   xor_2 : xor2_80 port map( a => s1, b => ci, o => s);
   and_1 : and2_81 port map( a => a, b => b, o => s2);
   and_2 : and2_80 port map( a => s1, b => ci, o => s3);
   or_1 : or2_40 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_39 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_39;

architecture SYN_Structural of fa_39 is

   component or2_39
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_78
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_79
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_78
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_79
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_79 port map( a => a, b => b, o => s1);
   xor_2 : xor2_78 port map( a => s1, b => ci, o => s);
   and_1 : and2_79 port map( a => a, b => b, o => s2);
   and_2 : and2_78 port map( a => s1, b => ci, o => s3);
   or_1 : or2_39 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_38 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_38;

architecture SYN_Structural of fa_38 is

   component or2_38
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_76
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_77
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_76
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_77
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_77 port map( a => a, b => b, o => s1);
   xor_2 : xor2_76 port map( a => s1, b => ci, o => s);
   and_1 : and2_77 port map( a => a, b => b, o => s2);
   and_2 : and2_76 port map( a => s1, b => ci, o => s3);
   or_1 : or2_38 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_37 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_37;

architecture SYN_Structural of fa_37 is

   component or2_37
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_74
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_75
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_74
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_75
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_75 port map( a => a, b => b, o => s1);
   xor_2 : xor2_74 port map( a => s1, b => ci, o => s);
   and_1 : and2_75 port map( a => a, b => b, o => s2);
   and_2 : and2_74 port map( a => s1, b => ci, o => s3);
   or_1 : or2_37 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_36 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_36;

architecture SYN_Structural of fa_36 is

   component or2_36
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_72
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_73
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_72
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_73
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_73 port map( a => a, b => b, o => s1);
   xor_2 : xor2_72 port map( a => s1, b => ci, o => s);
   and_1 : and2_73 port map( a => a, b => b, o => s2);
   and_2 : and2_72 port map( a => s1, b => ci, o => s3);
   or_1 : or2_36 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_35 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_35;

architecture SYN_Structural of fa_35 is

   component or2_35
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_70
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_71
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_70
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_71
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_71 port map( a => a, b => b, o => s1);
   xor_2 : xor2_70 port map( a => s1, b => ci, o => s);
   and_1 : and2_71 port map( a => a, b => b, o => s2);
   and_2 : and2_70 port map( a => s1, b => ci, o => s3);
   or_1 : or2_35 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_34 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_34;

architecture SYN_Structural of fa_34 is

   component or2_34
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_68
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_69
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_68
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_69
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_69 port map( a => a, b => b, o => s1);
   xor_2 : xor2_68 port map( a => s1, b => ci, o => s);
   and_1 : and2_69 port map( a => a, b => b, o => s2);
   and_2 : and2_68 port map( a => s1, b => ci, o => s3);
   or_1 : or2_34 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_33 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_33;

architecture SYN_Structural of fa_33 is

   component or2_33
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_66
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_67
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_66
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_67
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_67 port map( a => a, b => b, o => s1);
   xor_2 : xor2_66 port map( a => s1, b => ci, o => s);
   and_1 : and2_67 port map( a => a, b => b, o => s2);
   and_2 : and2_66 port map( a => s1, b => ci, o => s3);
   or_1 : or2_33 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_32 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_32;

architecture SYN_Structural of fa_32 is

   component or2_32
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_64
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_65
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_64
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_65
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_65 port map( a => a, b => b, o => s1);
   xor_2 : xor2_64 port map( a => s1, b => ci, o => s);
   and_1 : and2_65 port map( a => a, b => b, o => s2);
   and_2 : and2_64 port map( a => s1, b => ci, o => s3);
   or_1 : or2_32 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_31 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_31;

architecture SYN_Structural of fa_31 is

   component or2_31
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_61
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_62
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_61
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_62
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_62 port map( a => a, b => b, o => s1);
   xor_2 : xor2_61 port map( a => s1, b => ci, o => s);
   and_1 : and2_62 port map( a => a, b => b, o => s2);
   and_2 : and2_61 port map( a => s1, b => ci, o => s3);
   or_1 : or2_31 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_30 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_30;

architecture SYN_Structural of fa_30 is

   component or2_30
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_59
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_60
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_59
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_60
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_60 port map( a => a, b => b, o => s1);
   xor_2 : xor2_59 port map( a => s1, b => ci, o => s);
   and_1 : and2_60 port map( a => a, b => b, o => s2);
   and_2 : and2_59 port map( a => s1, b => ci, o => s3);
   or_1 : or2_30 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_29 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_29;

architecture SYN_Structural of fa_29 is

   component or2_29
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_57
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_58
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_57
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_58
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_58 port map( a => a, b => b, o => s1);
   xor_2 : xor2_57 port map( a => s1, b => ci, o => s);
   and_1 : and2_58 port map( a => a, b => b, o => s2);
   and_2 : and2_57 port map( a => s1, b => ci, o => s3);
   or_1 : or2_29 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_28 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_28;

architecture SYN_Structural of fa_28 is

   component or2_28
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_55
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_56
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_55
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_56
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_56 port map( a => a, b => b, o => s1);
   xor_2 : xor2_55 port map( a => s1, b => ci, o => s);
   and_1 : and2_56 port map( a => a, b => b, o => s2);
   and_2 : and2_55 port map( a => s1, b => ci, o => s3);
   or_1 : or2_28 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_27 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_27;

architecture SYN_Structural of fa_27 is

   component or2_27
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_53
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_54
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_53
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_54
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_54 port map( a => a, b => b, o => s1);
   xor_2 : xor2_53 port map( a => s1, b => ci, o => s);
   and_1 : and2_54 port map( a => a, b => b, o => s2);
   and_2 : and2_53 port map( a => s1, b => ci, o => s3);
   or_1 : or2_27 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_26 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_26;

architecture SYN_Structural of fa_26 is

   component or2_26
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_51
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_52
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_51
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_52
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_52 port map( a => a, b => b, o => s1);
   xor_2 : xor2_51 port map( a => s1, b => ci, o => s);
   and_1 : and2_52 port map( a => a, b => b, o => s2);
   and_2 : and2_51 port map( a => s1, b => ci, o => s3);
   or_1 : or2_26 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_25 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_25;

architecture SYN_Structural of fa_25 is

   component or2_25
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_49
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_50
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_49
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_50
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_50 port map( a => a, b => b, o => s1);
   xor_2 : xor2_49 port map( a => s1, b => ci, o => s);
   and_1 : and2_50 port map( a => a, b => b, o => s2);
   and_2 : and2_49 port map( a => s1, b => ci, o => s3);
   or_1 : or2_25 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_24 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_24;

architecture SYN_Structural of fa_24 is

   component or2_24
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_47
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_48
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_47
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_48
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_48 port map( a => a, b => b, o => s1);
   xor_2 : xor2_47 port map( a => s1, b => ci, o => s);
   and_1 : and2_48 port map( a => a, b => b, o => s2);
   and_2 : and2_47 port map( a => s1, b => ci, o => s3);
   or_1 : or2_24 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_23 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_23;

architecture SYN_Structural of fa_23 is

   component or2_23
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_45
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_46
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_45
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_46
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_46 port map( a => a, b => b, o => s1);
   xor_2 : xor2_45 port map( a => s1, b => ci, o => s);
   and_1 : and2_46 port map( a => a, b => b, o => s2);
   and_2 : and2_45 port map( a => s1, b => ci, o => s3);
   or_1 : or2_23 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_22 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_22;

architecture SYN_Structural of fa_22 is

   component or2_22
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_43
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_44
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_43
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_44
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_44 port map( a => a, b => b, o => s1);
   xor_2 : xor2_43 port map( a => s1, b => ci, o => s);
   and_1 : and2_44 port map( a => a, b => b, o => s2);
   and_2 : and2_43 port map( a => s1, b => ci, o => s3);
   or_1 : or2_22 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_21 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_21;

architecture SYN_Structural of fa_21 is

   component or2_21
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_41
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_42
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_41
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_42
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_42 port map( a => a, b => b, o => s1);
   xor_2 : xor2_41 port map( a => s1, b => ci, o => s);
   and_1 : and2_42 port map( a => a, b => b, o => s2);
   and_2 : and2_41 port map( a => s1, b => ci, o => s3);
   or_1 : or2_21 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_20 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_20;

architecture SYN_Structural of fa_20 is

   component or2_20
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_39
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_40
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_39
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_40
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_40 port map( a => a, b => b, o => s1);
   xor_2 : xor2_39 port map( a => s1, b => ci, o => s);
   and_1 : and2_40 port map( a => a, b => b, o => s2);
   and_2 : and2_39 port map( a => s1, b => ci, o => s3);
   or_1 : or2_20 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_19 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_19;

architecture SYN_Structural of fa_19 is

   component or2_19
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_37
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_38
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_37
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_38
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_38 port map( a => a, b => b, o => s1);
   xor_2 : xor2_37 port map( a => s1, b => ci, o => s);
   and_1 : and2_38 port map( a => a, b => b, o => s2);
   and_2 : and2_37 port map( a => s1, b => ci, o => s3);
   or_1 : or2_19 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_18 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_18;

architecture SYN_Structural of fa_18 is

   component or2_18
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_35
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_36
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_35
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_36
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_36 port map( a => a, b => b, o => s1);
   xor_2 : xor2_35 port map( a => s1, b => ci, o => s);
   and_1 : and2_36 port map( a => a, b => b, o => s2);
   and_2 : and2_35 port map( a => s1, b => ci, o => s3);
   or_1 : or2_18 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_17 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_17;

architecture SYN_Structural of fa_17 is

   component or2_17
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_33
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_34
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_33
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_34
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_34 port map( a => a, b => b, o => s1);
   xor_2 : xor2_33 port map( a => s1, b => ci, o => s);
   and_1 : and2_34 port map( a => a, b => b, o => s2);
   and_2 : and2_33 port map( a => s1, b => ci, o => s3);
   or_1 : or2_17 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_16 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_16;

architecture SYN_Structural of fa_16 is

   component or2_16
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_31
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_32
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_31
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_32
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_32 port map( a => a, b => b, o => s1);
   xor_2 : xor2_31 port map( a => s1, b => ci, o => s);
   and_1 : and2_32 port map( a => a, b => b, o => s2);
   and_2 : and2_31 port map( a => s1, b => ci, o => s3);
   or_1 : or2_16 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_15 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_15;

architecture SYN_Structural of fa_15 is

   component or2_15
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_29
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_30
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_29
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_30
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_30 port map( a => a, b => b, o => s1);
   xor_2 : xor2_29 port map( a => s1, b => ci, o => s);
   and_1 : and2_30 port map( a => a, b => b, o => s2);
   and_2 : and2_29 port map( a => s1, b => ci, o => s3);
   or_1 : or2_15 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_14 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_14;

architecture SYN_Structural of fa_14 is

   component or2_14
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_27
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_28
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_27
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_28
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_28 port map( a => a, b => b, o => s1);
   xor_2 : xor2_27 port map( a => s1, b => ci, o => s);
   and_1 : and2_28 port map( a => a, b => b, o => s2);
   and_2 : and2_27 port map( a => s1, b => ci, o => s3);
   or_1 : or2_14 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_13 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_13;

architecture SYN_Structural of fa_13 is

   component or2_13
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_25
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_26
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_25
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_26
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_26 port map( a => a, b => b, o => s1);
   xor_2 : xor2_25 port map( a => s1, b => ci, o => s);
   and_1 : and2_26 port map( a => a, b => b, o => s2);
   and_2 : and2_25 port map( a => s1, b => ci, o => s3);
   or_1 : or2_13 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_12 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_12;

architecture SYN_Structural of fa_12 is

   component or2_12
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_23
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_24
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_23
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_24
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_24 port map( a => a, b => b, o => s1);
   xor_2 : xor2_23 port map( a => s1, b => ci, o => s);
   and_1 : and2_24 port map( a => a, b => b, o => s2);
   and_2 : and2_23 port map( a => s1, b => ci, o => s3);
   or_1 : or2_12 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_11 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_11;

architecture SYN_Structural of fa_11 is

   component or2_11
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_21
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_22
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_21
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_22
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_22 port map( a => a, b => b, o => s1);
   xor_2 : xor2_21 port map( a => s1, b => ci, o => s);
   and_1 : and2_22 port map( a => a, b => b, o => s2);
   and_2 : and2_21 port map( a => s1, b => ci, o => s3);
   or_1 : or2_11 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_10 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_10;

architecture SYN_Structural of fa_10 is

   component or2_10
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_19
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_20
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_19
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_20
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_20 port map( a => a, b => b, o => s1);
   xor_2 : xor2_19 port map( a => s1, b => ci, o => s);
   and_1 : and2_20 port map( a => a, b => b, o => s2);
   and_2 : and2_19 port map( a => s1, b => ci, o => s3);
   or_1 : or2_10 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_9 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_9;

architecture SYN_Structural of fa_9 is

   component or2_9
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_17
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_18
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_17
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_18
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_18 port map( a => a, b => b, o => s1);
   xor_2 : xor2_17 port map( a => s1, b => ci, o => s);
   and_1 : and2_18 port map( a => a, b => b, o => s2);
   and_2 : and2_17 port map( a => s1, b => ci, o => s3);
   or_1 : or2_9 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_8 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_8;

architecture SYN_Structural of fa_8 is

   component or2_8
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_15
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_16
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_15
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_16
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_16 port map( a => a, b => b, o => s1);
   xor_2 : xor2_15 port map( a => s1, b => ci, o => s);
   and_1 : and2_16 port map( a => a, b => b, o => s2);
   and_2 : and2_15 port map( a => s1, b => ci, o => s3);
   or_1 : or2_8 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_7 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_7;

architecture SYN_Structural of fa_7 is

   component or2_7
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_13
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_14
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_13
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_14
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_14 port map( a => a, b => b, o => s1);
   xor_2 : xor2_13 port map( a => s1, b => ci, o => s);
   and_1 : and2_14 port map( a => a, b => b, o => s2);
   and_2 : and2_13 port map( a => s1, b => ci, o => s3);
   or_1 : or2_7 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_6 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_6;

architecture SYN_Structural of fa_6 is

   component or2_6
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_11
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_12
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_11
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_12
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_12 port map( a => a, b => b, o => s1);
   xor_2 : xor2_11 port map( a => s1, b => ci, o => s);
   and_1 : and2_12 port map( a => a, b => b, o => s2);
   and_2 : and2_11 port map( a => s1, b => ci, o => s3);
   or_1 : or2_6 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_5 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_5;

architecture SYN_Structural of fa_5 is

   component or2_5
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_9
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_10
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_9
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_10
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_10 port map( a => a, b => b, o => s1);
   xor_2 : xor2_9 port map( a => s1, b => ci, o => s);
   and_1 : and2_10 port map( a => a, b => b, o => s2);
   and_2 : and2_9 port map( a => s1, b => ci, o => s3);
   or_1 : or2_5 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_4 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_4;

architecture SYN_Structural of fa_4 is

   component or2_4
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_7
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_8
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_7
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_8
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_8 port map( a => a, b => b, o => s1);
   xor_2 : xor2_7 port map( a => s1, b => ci, o => s);
   and_1 : and2_8 port map( a => a, b => b, o => s2);
   and_2 : and2_7 port map( a => s1, b => ci, o => s3);
   or_1 : or2_4 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_3 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_3;

architecture SYN_Structural of fa_3 is

   component or2_3
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_5
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_6
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_5
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_6
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_6 port map( a => a, b => b, o => s1);
   xor_2 : xor2_5 port map( a => s1, b => ci, o => s);
   and_1 : and2_6 port map( a => a, b => b, o => s2);
   and_2 : and2_5 port map( a => s1, b => ci, o => s3);
   or_1 : or2_3 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_2 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_2;

architecture SYN_Structural of fa_2 is

   component or2_2
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_3
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_4
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_3
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_4
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_4 port map( a => a, b => b, o => s1);
   xor_2 : xor2_3 port map( a => s1, b => ci, o => s);
   and_1 : and2_4 port map( a => a, b => b, o => s2);
   and_2 : and2_3 port map( a => s1, b => ci, o => s3);
   or_1 : or2_2 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_1 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_1;

architecture SYN_Structural of fa_1 is

   component or2_1
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_1
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_2
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_1
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_2
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_2 port map( a => a, b => b, o => s1);
   xor_2 : xor2_1 port map( a => s1, b => ci, o => s);
   and_1 : and2_2 port map( a => a, b => b, o => s2);
   and_2 : and2_1 port map( a => s1, b => ci, o => s3);
   or_1 : or2_1 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity half_adder_6 is

   port( a, b : in std_logic;  co, s : out std_logic);

end half_adder_6;

architecture SYN_Structural of half_adder_6 is

   component xor2_378
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_378
      port( a, b : in std_logic;  o : out std_logic);
   end component;

begin
   
   carry : and2_378 port map( a => a, b => b, o => co);
   sum : xor2_378 port map( a => a, b => b, o => s);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity half_adder_5 is

   port( a, b : in std_logic;  co, s : out std_logic);

end half_adder_5;

architecture SYN_Structural of half_adder_5 is

   component xor2_315
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_315
      port( a, b : in std_logic;  o : out std_logic);
   end component;

begin
   
   carry : and2_315 port map( a => a, b => b, o => co);
   sum : xor2_315 port map( a => a, b => b, o => s);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity half_adder_4 is

   port( a, b : in std_logic;  co, s : out std_logic);

end half_adder_4;

architecture SYN_Structural of half_adder_4 is

   component xor2_252
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_252
      port( a, b : in std_logic;  o : out std_logic);
   end component;

begin
   
   carry : and2_252 port map( a => a, b => b, o => co);
   sum : xor2_252 port map( a => a, b => b, o => s);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity half_adder_3 is

   port( a, b : in std_logic;  co, s : out std_logic);

end half_adder_3;

architecture SYN_Structural of half_adder_3 is

   component xor2_189
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_189
      port( a, b : in std_logic;  o : out std_logic);
   end component;

begin
   
   carry : and2_189 port map( a => a, b => b, o => co);
   sum : xor2_189 port map( a => a, b => b, o => s);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity half_adder_2 is

   port( a, b : in std_logic;  co, s : out std_logic);

end half_adder_2;

architecture SYN_Structural of half_adder_2 is

   component xor2_126
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_126
      port( a, b : in std_logic;  o : out std_logic);
   end component;

begin
   
   carry : and2_126 port map( a => a, b => b, o => co);
   sum : xor2_126 port map( a => a, b => b, o => s);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity half_adder_1 is

   port( a, b : in std_logic;  co, s : out std_logic);

end half_adder_1;

architecture SYN_Structural of half_adder_1 is

   component xor2_63
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_63
      port( a, b : in std_logic;  o : out std_logic);
   end component;

begin
   
   carry : and2_63 port map( a => a, b => b, o => co);
   sum : xor2_63 port map( a => a, b => b, o => s);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_15 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_15;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_57
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_58
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_59
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_60
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_60 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_59 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_58 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_57 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_14 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_14;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_53
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_54
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_55
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_56
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_56 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_55 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_54 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_53 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_13 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_13;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_49
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_50
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_51
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_52
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_52 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_51 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_50 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_49 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_12 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_12;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_45
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_46
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_47
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_48
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_48 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_47 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_46 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_45 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_11 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_11;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_41
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_42
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_43
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_44
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_44 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_43 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_42 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_41 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_10 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_10;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_37
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_38
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_39
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_40
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_40 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_39 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_38 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_37 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_9 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_9;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_33
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_34
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_35
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_36
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_36 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_35 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_34 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_33 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_8 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_8;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_29
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_30
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_31
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_32
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_32 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_31 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_30 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_29 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_7 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_7;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_25
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_26
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_27
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_28
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_28 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_27 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_26 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_25 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_6 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_6;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_21
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_22
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_23
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_24
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_24 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_23 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_22 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_21 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_5 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_5;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_17
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_18
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_19
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_20
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_20 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_19 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_18 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_17 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_4 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_4;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_13
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_14
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_15
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_16
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_16 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_15 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_14 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_13 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_3 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_3;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_9
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_10
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_11
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_12
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_12 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_11 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_10 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_9 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_2 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_2;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_5
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_6
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_7
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_8
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_8 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_7 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_6 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_5 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_1 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_1;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_1
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_2
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_3
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_4
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_4 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_3 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_2 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_1 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_7 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_7;

architecture SYN_specification of g_block_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_6 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_6;

architecture SYN_specification of g_block_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_5 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_5;

architecture SYN_specification of g_block_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_4 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_4;

architecture SYN_specification of g_block_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_3 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_3;

architecture SYN_specification of g_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_2 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_2;

architecture SYN_specification of g_block_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_1 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_1;

architecture SYN_specification of g_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_26 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_26;

architecture SYN_specification of pg_block_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_25 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_25;

architecture SYN_specification of pg_block_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_24 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_24;

architecture SYN_specification of pg_block_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_23 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_23;

architecture SYN_specification of pg_block_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_22 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_22;

architecture SYN_specification of pg_block_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_21 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_21;

architecture SYN_specification of pg_block_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_20 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_20;

architecture SYN_specification of pg_block_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_19 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_19;

architecture SYN_specification of pg_block_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_18 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_18;

architecture SYN_specification of pg_block_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_17 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_17;

architecture SYN_specification of pg_block_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_16 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_16;

architecture SYN_specification of pg_block_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_15 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_15;

architecture SYN_specification of pg_block_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_14 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_14;

architecture SYN_specification of pg_block_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_13 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_13;

architecture SYN_specification of pg_block_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_12 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_12;

architecture SYN_specification of pg_block_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_11 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_11;

architecture SYN_specification of pg_block_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_10 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_10;

architecture SYN_specification of pg_block_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_9 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_9;

architecture SYN_specification of pg_block_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_8 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_8;

architecture SYN_specification of pg_block_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_7 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_7;

architecture SYN_specification of pg_block_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_6 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_6;

architecture SYN_specification of pg_block_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_5 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_5;

architecture SYN_specification of pg_block_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_4 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_4;

architecture SYN_specification of pg_block_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_3 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_3;

architecture SYN_specification of pg_block_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_2 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_2;

architecture SYN_specification of pg_block_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_1 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_1;

architecture SYN_specification of pg_block_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N40_3 is

   port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (39 downto 0));

end MUX21_N40_3;

architecture SYN_beh of MUX21_N40_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));
   U2 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U3 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U4 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U5 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U6 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U7 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U8 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U9 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U10 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U11 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U12 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U13 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U14 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U15 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U16 : MUX2_X1 port map( A => a(39), B => b(39), S => sel, Z => y(39));
   U17 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U18 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U19 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U20 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U21 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U22 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U23 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U24 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U25 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U26 : MUX2_X1 port map( A => a(32), B => b(32), S => sel, Z => y(32));
   U27 : MUX2_X1 port map( A => a(33), B => b(33), S => sel, Z => y(33));
   U28 : MUX2_X1 port map( A => a(34), B => b(34), S => sel, Z => y(34));
   U29 : MUX2_X1 port map( A => a(35), B => b(35), S => sel, Z => y(35));
   U30 : MUX2_X1 port map( A => a(36), B => b(36), S => sel, Z => y(36));
   U31 : MUX2_X1 port map( A => a(37), B => b(37), S => sel, Z => y(37));
   U32 : MUX2_X1 port map( A => a(38), B => b(38), S => sel, Z => y(38));
   U33 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U34 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U35 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U36 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U37 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U38 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U39 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U40 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N40_2 is

   port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (39 downto 0));

end MUX21_N40_2;

architecture SYN_beh of MUX21_N40_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));
   U2 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U3 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U4 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U5 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U6 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U7 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U8 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U9 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U10 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U11 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U12 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U13 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U14 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U15 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U16 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U17 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U18 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U19 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U20 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U21 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U22 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U23 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U24 : MUX2_X1 port map( A => a(39), B => b(39), S => sel, Z => y(39));
   U25 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U26 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U27 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U28 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U29 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U30 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U31 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U32 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U33 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U34 : MUX2_X1 port map( A => a(32), B => b(32), S => sel, Z => y(32));
   U35 : MUX2_X1 port map( A => a(33), B => b(33), S => sel, Z => y(33));
   U36 : MUX2_X1 port map( A => a(34), B => b(34), S => sel, Z => y(34));
   U37 : MUX2_X1 port map( A => a(35), B => b(35), S => sel, Z => y(35));
   U38 : MUX2_X1 port map( A => a(36), B => b(36), S => sel, Z => y(36));
   U39 : MUX2_X1 port map( A => a(37), B => b(37), S => sel, Z => y(37));
   U40 : MUX2_X1 port map( A => a(38), B => b(38), S => sel, Z => y(38));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N40_1 is

   port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (39 downto 0));

end MUX21_N40_1;

architecture SYN_beh of MUX21_N40_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));
   U2 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U3 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U4 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U5 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U6 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U7 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U8 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U9 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U10 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U11 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U12 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U13 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U14 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U15 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U16 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U17 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U18 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U19 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U20 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U21 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U22 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U23 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U24 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U25 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U26 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U27 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U28 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U29 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U30 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U31 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U32 : MUX2_X1 port map( A => a(39), B => b(39), S => sel, Z => y(39));
   U33 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U34 : MUX2_X1 port map( A => a(32), B => b(32), S => sel, Z => y(32));
   U35 : MUX2_X1 port map( A => a(33), B => b(33), S => sel, Z => y(33));
   U36 : MUX2_X1 port map( A => a(34), B => b(34), S => sel, Z => y(34));
   U37 : MUX2_X1 port map( A => a(35), B => b(35), S => sel, Z => y(35));
   U38 : MUX2_X1 port map( A => a(36), B => b(36), S => sel, Z => y(36));
   U39 : MUX2_X1 port map( A => a(37), B => b(37), S => sel, Z => y(37));
   U40 : MUX2_X1 port map( A => a(38), B => b(38), S => sel, Z => y(38));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity rca_signed_NBIT32_6 is

   port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : out
         std_logic_vector (31 downto 0));

end rca_signed_NBIT32_6;

architecture SYN_Structural of rca_signed_NBIT32_6 is

   component fa_156
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_157
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_158
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_159
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_160
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_161
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_162
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_163
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_164
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_165
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_166
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_167
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_168
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_169
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_170
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_171
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_172
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_173
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_174
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_175
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_176
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_177
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_178
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_179
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_180
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_181
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_182
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_183
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_184
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_185
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_186
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component half_adder_6
      port( a, b : in std_logic;  co, s : out std_logic);
   end component;
   
   signal carry_s_30_port, carry_s_29_port, carry_s_28_port, carry_s_27_port, 
      carry_s_26_port, carry_s_25_port, carry_s_24_port, carry_s_23_port, 
      carry_s_22_port, carry_s_21_port, carry_s_20_port, carry_s_19_port, 
      carry_s_18_port, carry_s_17_port, carry_s_16_port, carry_s_15_port, 
      carry_s_14_port, carry_s_13_port, carry_s_12_port, carry_s_11_port, 
      carry_s_10_port, carry_s_9_port, carry_s_8_port, carry_s_7_port, 
      carry_s_6_port, carry_s_5_port, carry_s_4_port, carry_s_3_port, 
      carry_s_2_port, carry_s_1_port, carry_s_0_port : std_logic;

begin
   
   ha : half_adder_6 port map( a => a(0), b => b(0), co => carry_s_0_port, s =>
                           s(0));
   fa_i_1 : fa_186 port map( a => a(1), b => b(1), ci => carry_s_0_port, co => 
                           carry_s_1_port, s => s(1));
   fa_i_2 : fa_185 port map( a => a(2), b => b(2), ci => carry_s_1_port, co => 
                           carry_s_2_port, s => s(2));
   fa_i_3 : fa_184 port map( a => a(3), b => b(3), ci => carry_s_2_port, co => 
                           carry_s_3_port, s => s(3));
   fa_i_4 : fa_183 port map( a => a(4), b => b(4), ci => carry_s_3_port, co => 
                           carry_s_4_port, s => s(4));
   fa_i_5 : fa_182 port map( a => a(5), b => b(5), ci => carry_s_4_port, co => 
                           carry_s_5_port, s => s(5));
   fa_i_6 : fa_181 port map( a => a(6), b => b(6), ci => carry_s_5_port, co => 
                           carry_s_6_port, s => s(6));
   fa_i_7 : fa_180 port map( a => a(7), b => b(7), ci => carry_s_6_port, co => 
                           carry_s_7_port, s => s(7));
   fa_i_8 : fa_179 port map( a => a(8), b => b(8), ci => carry_s_7_port, co => 
                           carry_s_8_port, s => s(8));
   fa_i_9 : fa_178 port map( a => a(9), b => b(9), ci => carry_s_8_port, co => 
                           carry_s_9_port, s => s(9));
   fa_i_10 : fa_177 port map( a => a(10), b => b(10), ci => carry_s_9_port, co 
                           => carry_s_10_port, s => s(10));
   fa_i_11 : fa_176 port map( a => a(11), b => b(11), ci => carry_s_10_port, co
                           => carry_s_11_port, s => s(11));
   fa_i_12 : fa_175 port map( a => a(12), b => b(12), ci => carry_s_11_port, co
                           => carry_s_12_port, s => s(12));
   fa_i_13 : fa_174 port map( a => a(13), b => b(13), ci => carry_s_12_port, co
                           => carry_s_13_port, s => s(13));
   fa_i_14 : fa_173 port map( a => a(14), b => b(14), ci => carry_s_13_port, co
                           => carry_s_14_port, s => s(14));
   fa_i_15 : fa_172 port map( a => a(15), b => b(15), ci => carry_s_14_port, co
                           => carry_s_15_port, s => s(15));
   fa_i_16 : fa_171 port map( a => a(16), b => b(16), ci => carry_s_15_port, co
                           => carry_s_16_port, s => s(16));
   fa_i_17 : fa_170 port map( a => a(17), b => b(17), ci => carry_s_16_port, co
                           => carry_s_17_port, s => s(17));
   fa_i_18 : fa_169 port map( a => a(18), b => b(18), ci => carry_s_17_port, co
                           => carry_s_18_port, s => s(18));
   fa_i_19 : fa_168 port map( a => a(19), b => b(19), ci => carry_s_18_port, co
                           => carry_s_19_port, s => s(19));
   fa_i_20 : fa_167 port map( a => a(20), b => b(20), ci => carry_s_19_port, co
                           => carry_s_20_port, s => s(20));
   fa_i_21 : fa_166 port map( a => a(21), b => b(21), ci => carry_s_20_port, co
                           => carry_s_21_port, s => s(21));
   fa_i_22 : fa_165 port map( a => a(22), b => b(22), ci => carry_s_21_port, co
                           => carry_s_22_port, s => s(22));
   fa_i_23 : fa_164 port map( a => a(23), b => b(23), ci => carry_s_22_port, co
                           => carry_s_23_port, s => s(23));
   fa_i_24 : fa_163 port map( a => a(24), b => b(24), ci => carry_s_23_port, co
                           => carry_s_24_port, s => s(24));
   fa_i_25 : fa_162 port map( a => a(25), b => b(25), ci => carry_s_24_port, co
                           => carry_s_25_port, s => s(25));
   fa_i_26 : fa_161 port map( a => a(26), b => b(26), ci => carry_s_25_port, co
                           => carry_s_26_port, s => s(26));
   fa_i_27 : fa_160 port map( a => a(27), b => b(27), ci => carry_s_26_port, co
                           => carry_s_27_port, s => s(27));
   fa_i_28 : fa_159 port map( a => a(28), b => b(28), ci => carry_s_27_port, co
                           => carry_s_28_port, s => s(28));
   fa_i_29 : fa_158 port map( a => a(29), b => b(29), ci => carry_s_28_port, co
                           => carry_s_29_port, s => s(29));
   fa_i_30 : fa_157 port map( a => a(30), b => b(30), ci => carry_s_29_port, co
                           => carry_s_30_port, s => s(30));
   fa_i_31 : fa_156 port map( a => a(31), b => b(31), ci => carry_s_30_port, co
                           => c, s => s(31));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity rca_signed_NBIT32_5 is

   port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : out
         std_logic_vector (31 downto 0));

end rca_signed_NBIT32_5;

architecture SYN_Structural of rca_signed_NBIT32_5 is

   component fa_125
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_126
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_127
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_128
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_129
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_130
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_131
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_132
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_133
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_134
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_135
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_136
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_137
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_138
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_139
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_140
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_141
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_142
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_143
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_144
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_145
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_146
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_147
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_148
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_149
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_150
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_151
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_152
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_153
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_154
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_155
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component half_adder_5
      port( a, b : in std_logic;  co, s : out std_logic);
   end component;
   
   signal carry_s_30_port, carry_s_29_port, carry_s_28_port, carry_s_27_port, 
      carry_s_26_port, carry_s_25_port, carry_s_24_port, carry_s_23_port, 
      carry_s_22_port, carry_s_21_port, carry_s_20_port, carry_s_19_port, 
      carry_s_18_port, carry_s_17_port, carry_s_16_port, carry_s_15_port, 
      carry_s_14_port, carry_s_13_port, carry_s_12_port, carry_s_11_port, 
      carry_s_10_port, carry_s_9_port, carry_s_8_port, carry_s_7_port, 
      carry_s_6_port, carry_s_5_port, carry_s_4_port, carry_s_3_port, 
      carry_s_2_port, carry_s_1_port, carry_s_0_port : std_logic;

begin
   
   ha : half_adder_5 port map( a => a(0), b => b(0), co => carry_s_0_port, s =>
                           s(0));
   fa_i_1 : fa_155 port map( a => a(1), b => b(1), ci => carry_s_0_port, co => 
                           carry_s_1_port, s => s(1));
   fa_i_2 : fa_154 port map( a => a(2), b => b(2), ci => carry_s_1_port, co => 
                           carry_s_2_port, s => s(2));
   fa_i_3 : fa_153 port map( a => a(3), b => b(3), ci => carry_s_2_port, co => 
                           carry_s_3_port, s => s(3));
   fa_i_4 : fa_152 port map( a => a(4), b => b(4), ci => carry_s_3_port, co => 
                           carry_s_4_port, s => s(4));
   fa_i_5 : fa_151 port map( a => a(5), b => b(5), ci => carry_s_4_port, co => 
                           carry_s_5_port, s => s(5));
   fa_i_6 : fa_150 port map( a => a(6), b => b(6), ci => carry_s_5_port, co => 
                           carry_s_6_port, s => s(6));
   fa_i_7 : fa_149 port map( a => a(7), b => b(7), ci => carry_s_6_port, co => 
                           carry_s_7_port, s => s(7));
   fa_i_8 : fa_148 port map( a => a(8), b => b(8), ci => carry_s_7_port, co => 
                           carry_s_8_port, s => s(8));
   fa_i_9 : fa_147 port map( a => a(9), b => b(9), ci => carry_s_8_port, co => 
                           carry_s_9_port, s => s(9));
   fa_i_10 : fa_146 port map( a => a(10), b => b(10), ci => carry_s_9_port, co 
                           => carry_s_10_port, s => s(10));
   fa_i_11 : fa_145 port map( a => a(11), b => b(11), ci => carry_s_10_port, co
                           => carry_s_11_port, s => s(11));
   fa_i_12 : fa_144 port map( a => a(12), b => b(12), ci => carry_s_11_port, co
                           => carry_s_12_port, s => s(12));
   fa_i_13 : fa_143 port map( a => a(13), b => b(13), ci => carry_s_12_port, co
                           => carry_s_13_port, s => s(13));
   fa_i_14 : fa_142 port map( a => a(14), b => b(14), ci => carry_s_13_port, co
                           => carry_s_14_port, s => s(14));
   fa_i_15 : fa_141 port map( a => a(15), b => b(15), ci => carry_s_14_port, co
                           => carry_s_15_port, s => s(15));
   fa_i_16 : fa_140 port map( a => a(16), b => b(16), ci => carry_s_15_port, co
                           => carry_s_16_port, s => s(16));
   fa_i_17 : fa_139 port map( a => a(17), b => b(17), ci => carry_s_16_port, co
                           => carry_s_17_port, s => s(17));
   fa_i_18 : fa_138 port map( a => a(18), b => b(18), ci => carry_s_17_port, co
                           => carry_s_18_port, s => s(18));
   fa_i_19 : fa_137 port map( a => a(19), b => b(19), ci => carry_s_18_port, co
                           => carry_s_19_port, s => s(19));
   fa_i_20 : fa_136 port map( a => a(20), b => b(20), ci => carry_s_19_port, co
                           => carry_s_20_port, s => s(20));
   fa_i_21 : fa_135 port map( a => a(21), b => b(21), ci => carry_s_20_port, co
                           => carry_s_21_port, s => s(21));
   fa_i_22 : fa_134 port map( a => a(22), b => b(22), ci => carry_s_21_port, co
                           => carry_s_22_port, s => s(22));
   fa_i_23 : fa_133 port map( a => a(23), b => b(23), ci => carry_s_22_port, co
                           => carry_s_23_port, s => s(23));
   fa_i_24 : fa_132 port map( a => a(24), b => b(24), ci => carry_s_23_port, co
                           => carry_s_24_port, s => s(24));
   fa_i_25 : fa_131 port map( a => a(25), b => b(25), ci => carry_s_24_port, co
                           => carry_s_25_port, s => s(25));
   fa_i_26 : fa_130 port map( a => a(26), b => b(26), ci => carry_s_25_port, co
                           => carry_s_26_port, s => s(26));
   fa_i_27 : fa_129 port map( a => a(27), b => b(27), ci => carry_s_26_port, co
                           => carry_s_27_port, s => s(27));
   fa_i_28 : fa_128 port map( a => a(28), b => b(28), ci => carry_s_27_port, co
                           => carry_s_28_port, s => s(28));
   fa_i_29 : fa_127 port map( a => a(29), b => b(29), ci => carry_s_28_port, co
                           => carry_s_29_port, s => s(29));
   fa_i_30 : fa_126 port map( a => a(30), b => b(30), ci => carry_s_29_port, co
                           => carry_s_30_port, s => s(30));
   fa_i_31 : fa_125 port map( a => a(31), b => b(31), ci => carry_s_30_port, co
                           => c, s => s(31));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity rca_signed_NBIT32_4 is

   port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : out
         std_logic_vector (31 downto 0));

end rca_signed_NBIT32_4;

architecture SYN_Structural of rca_signed_NBIT32_4 is

   component fa_94
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_95
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_96
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_97
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_98
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_99
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_100
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_101
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_102
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_103
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_104
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_105
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_106
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_107
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_108
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_109
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_110
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_111
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_112
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_113
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_114
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_115
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_116
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_117
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_118
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_119
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_120
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_121
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_122
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_123
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_124
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component half_adder_4
      port( a, b : in std_logic;  co, s : out std_logic);
   end component;
   
   signal carry_s_30_port, carry_s_29_port, carry_s_28_port, carry_s_27_port, 
      carry_s_26_port, carry_s_25_port, carry_s_24_port, carry_s_23_port, 
      carry_s_22_port, carry_s_21_port, carry_s_20_port, carry_s_19_port, 
      carry_s_18_port, carry_s_17_port, carry_s_16_port, carry_s_15_port, 
      carry_s_14_port, carry_s_13_port, carry_s_12_port, carry_s_11_port, 
      carry_s_10_port, carry_s_9_port, carry_s_8_port, carry_s_7_port, 
      carry_s_6_port, carry_s_5_port, carry_s_4_port, carry_s_3_port, 
      carry_s_2_port, carry_s_1_port, carry_s_0_port : std_logic;

begin
   
   ha : half_adder_4 port map( a => a(0), b => b(0), co => carry_s_0_port, s =>
                           s(0));
   fa_i_1 : fa_124 port map( a => a(1), b => b(1), ci => carry_s_0_port, co => 
                           carry_s_1_port, s => s(1));
   fa_i_2 : fa_123 port map( a => a(2), b => b(2), ci => carry_s_1_port, co => 
                           carry_s_2_port, s => s(2));
   fa_i_3 : fa_122 port map( a => a(3), b => b(3), ci => carry_s_2_port, co => 
                           carry_s_3_port, s => s(3));
   fa_i_4 : fa_121 port map( a => a(4), b => b(4), ci => carry_s_3_port, co => 
                           carry_s_4_port, s => s(4));
   fa_i_5 : fa_120 port map( a => a(5), b => b(5), ci => carry_s_4_port, co => 
                           carry_s_5_port, s => s(5));
   fa_i_6 : fa_119 port map( a => a(6), b => b(6), ci => carry_s_5_port, co => 
                           carry_s_6_port, s => s(6));
   fa_i_7 : fa_118 port map( a => a(7), b => b(7), ci => carry_s_6_port, co => 
                           carry_s_7_port, s => s(7));
   fa_i_8 : fa_117 port map( a => a(8), b => b(8), ci => carry_s_7_port, co => 
                           carry_s_8_port, s => s(8));
   fa_i_9 : fa_116 port map( a => a(9), b => b(9), ci => carry_s_8_port, co => 
                           carry_s_9_port, s => s(9));
   fa_i_10 : fa_115 port map( a => a(10), b => b(10), ci => carry_s_9_port, co 
                           => carry_s_10_port, s => s(10));
   fa_i_11 : fa_114 port map( a => a(11), b => b(11), ci => carry_s_10_port, co
                           => carry_s_11_port, s => s(11));
   fa_i_12 : fa_113 port map( a => a(12), b => b(12), ci => carry_s_11_port, co
                           => carry_s_12_port, s => s(12));
   fa_i_13 : fa_112 port map( a => a(13), b => b(13), ci => carry_s_12_port, co
                           => carry_s_13_port, s => s(13));
   fa_i_14 : fa_111 port map( a => a(14), b => b(14), ci => carry_s_13_port, co
                           => carry_s_14_port, s => s(14));
   fa_i_15 : fa_110 port map( a => a(15), b => b(15), ci => carry_s_14_port, co
                           => carry_s_15_port, s => s(15));
   fa_i_16 : fa_109 port map( a => a(16), b => b(16), ci => carry_s_15_port, co
                           => carry_s_16_port, s => s(16));
   fa_i_17 : fa_108 port map( a => a(17), b => b(17), ci => carry_s_16_port, co
                           => carry_s_17_port, s => s(17));
   fa_i_18 : fa_107 port map( a => a(18), b => b(18), ci => carry_s_17_port, co
                           => carry_s_18_port, s => s(18));
   fa_i_19 : fa_106 port map( a => a(19), b => b(19), ci => carry_s_18_port, co
                           => carry_s_19_port, s => s(19));
   fa_i_20 : fa_105 port map( a => a(20), b => b(20), ci => carry_s_19_port, co
                           => carry_s_20_port, s => s(20));
   fa_i_21 : fa_104 port map( a => a(21), b => b(21), ci => carry_s_20_port, co
                           => carry_s_21_port, s => s(21));
   fa_i_22 : fa_103 port map( a => a(22), b => b(22), ci => carry_s_21_port, co
                           => carry_s_22_port, s => s(22));
   fa_i_23 : fa_102 port map( a => a(23), b => b(23), ci => carry_s_22_port, co
                           => carry_s_23_port, s => s(23));
   fa_i_24 : fa_101 port map( a => a(24), b => b(24), ci => carry_s_23_port, co
                           => carry_s_24_port, s => s(24));
   fa_i_25 : fa_100 port map( a => a(25), b => b(25), ci => carry_s_24_port, co
                           => carry_s_25_port, s => s(25));
   fa_i_26 : fa_99 port map( a => a(26), b => b(26), ci => carry_s_25_port, co 
                           => carry_s_26_port, s => s(26));
   fa_i_27 : fa_98 port map( a => a(27), b => b(27), ci => carry_s_26_port, co 
                           => carry_s_27_port, s => s(27));
   fa_i_28 : fa_97 port map( a => a(28), b => b(28), ci => carry_s_27_port, co 
                           => carry_s_28_port, s => s(28));
   fa_i_29 : fa_96 port map( a => a(29), b => b(29), ci => carry_s_28_port, co 
                           => carry_s_29_port, s => s(29));
   fa_i_30 : fa_95 port map( a => a(30), b => b(30), ci => carry_s_29_port, co 
                           => carry_s_30_port, s => s(30));
   fa_i_31 : fa_94 port map( a => a(31), b => b(31), ci => carry_s_30_port, co 
                           => c, s => s(31));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity rca_signed_NBIT32_3 is

   port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : out
         std_logic_vector (31 downto 0));

end rca_signed_NBIT32_3;

architecture SYN_Structural of rca_signed_NBIT32_3 is

   component fa_63
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_64
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_65
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_66
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_67
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_68
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_69
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_70
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_71
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_72
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_73
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_74
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_75
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_76
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_77
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_78
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_79
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_80
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_81
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_82
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_83
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_84
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_85
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_86
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_87
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_88
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_89
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_90
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_91
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_92
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_93
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component half_adder_3
      port( a, b : in std_logic;  co, s : out std_logic);
   end component;
   
   signal carry_s_30_port, carry_s_29_port, carry_s_28_port, carry_s_27_port, 
      carry_s_26_port, carry_s_25_port, carry_s_24_port, carry_s_23_port, 
      carry_s_22_port, carry_s_21_port, carry_s_20_port, carry_s_19_port, 
      carry_s_18_port, carry_s_17_port, carry_s_16_port, carry_s_15_port, 
      carry_s_14_port, carry_s_13_port, carry_s_12_port, carry_s_11_port, 
      carry_s_10_port, carry_s_9_port, carry_s_8_port, carry_s_7_port, 
      carry_s_6_port, carry_s_5_port, carry_s_4_port, carry_s_3_port, 
      carry_s_2_port, carry_s_1_port, carry_s_0_port : std_logic;

begin
   
   ha : half_adder_3 port map( a => a(0), b => b(0), co => carry_s_0_port, s =>
                           s(0));
   fa_i_1 : fa_93 port map( a => a(1), b => b(1), ci => carry_s_0_port, co => 
                           carry_s_1_port, s => s(1));
   fa_i_2 : fa_92 port map( a => a(2), b => b(2), ci => carry_s_1_port, co => 
                           carry_s_2_port, s => s(2));
   fa_i_3 : fa_91 port map( a => a(3), b => b(3), ci => carry_s_2_port, co => 
                           carry_s_3_port, s => s(3));
   fa_i_4 : fa_90 port map( a => a(4), b => b(4), ci => carry_s_3_port, co => 
                           carry_s_4_port, s => s(4));
   fa_i_5 : fa_89 port map( a => a(5), b => b(5), ci => carry_s_4_port, co => 
                           carry_s_5_port, s => s(5));
   fa_i_6 : fa_88 port map( a => a(6), b => b(6), ci => carry_s_5_port, co => 
                           carry_s_6_port, s => s(6));
   fa_i_7 : fa_87 port map( a => a(7), b => b(7), ci => carry_s_6_port, co => 
                           carry_s_7_port, s => s(7));
   fa_i_8 : fa_86 port map( a => a(8), b => b(8), ci => carry_s_7_port, co => 
                           carry_s_8_port, s => s(8));
   fa_i_9 : fa_85 port map( a => a(9), b => b(9), ci => carry_s_8_port, co => 
                           carry_s_9_port, s => s(9));
   fa_i_10 : fa_84 port map( a => a(10), b => b(10), ci => carry_s_9_port, co 
                           => carry_s_10_port, s => s(10));
   fa_i_11 : fa_83 port map( a => a(11), b => b(11), ci => carry_s_10_port, co 
                           => carry_s_11_port, s => s(11));
   fa_i_12 : fa_82 port map( a => a(12), b => b(12), ci => carry_s_11_port, co 
                           => carry_s_12_port, s => s(12));
   fa_i_13 : fa_81 port map( a => a(13), b => b(13), ci => carry_s_12_port, co 
                           => carry_s_13_port, s => s(13));
   fa_i_14 : fa_80 port map( a => a(14), b => b(14), ci => carry_s_13_port, co 
                           => carry_s_14_port, s => s(14));
   fa_i_15 : fa_79 port map( a => a(15), b => b(15), ci => carry_s_14_port, co 
                           => carry_s_15_port, s => s(15));
   fa_i_16 : fa_78 port map( a => a(16), b => b(16), ci => carry_s_15_port, co 
                           => carry_s_16_port, s => s(16));
   fa_i_17 : fa_77 port map( a => a(17), b => b(17), ci => carry_s_16_port, co 
                           => carry_s_17_port, s => s(17));
   fa_i_18 : fa_76 port map( a => a(18), b => b(18), ci => carry_s_17_port, co 
                           => carry_s_18_port, s => s(18));
   fa_i_19 : fa_75 port map( a => a(19), b => b(19), ci => carry_s_18_port, co 
                           => carry_s_19_port, s => s(19));
   fa_i_20 : fa_74 port map( a => a(20), b => b(20), ci => carry_s_19_port, co 
                           => carry_s_20_port, s => s(20));
   fa_i_21 : fa_73 port map( a => a(21), b => b(21), ci => carry_s_20_port, co 
                           => carry_s_21_port, s => s(21));
   fa_i_22 : fa_72 port map( a => a(22), b => b(22), ci => carry_s_21_port, co 
                           => carry_s_22_port, s => s(22));
   fa_i_23 : fa_71 port map( a => a(23), b => b(23), ci => carry_s_22_port, co 
                           => carry_s_23_port, s => s(23));
   fa_i_24 : fa_70 port map( a => a(24), b => b(24), ci => carry_s_23_port, co 
                           => carry_s_24_port, s => s(24));
   fa_i_25 : fa_69 port map( a => a(25), b => b(25), ci => carry_s_24_port, co 
                           => carry_s_25_port, s => s(25));
   fa_i_26 : fa_68 port map( a => a(26), b => b(26), ci => carry_s_25_port, co 
                           => carry_s_26_port, s => s(26));
   fa_i_27 : fa_67 port map( a => a(27), b => b(27), ci => carry_s_26_port, co 
                           => carry_s_27_port, s => s(27));
   fa_i_28 : fa_66 port map( a => a(28), b => b(28), ci => carry_s_27_port, co 
                           => carry_s_28_port, s => s(28));
   fa_i_29 : fa_65 port map( a => a(29), b => b(29), ci => carry_s_28_port, co 
                           => carry_s_29_port, s => s(29));
   fa_i_30 : fa_64 port map( a => a(30), b => b(30), ci => carry_s_29_port, co 
                           => carry_s_30_port, s => s(30));
   fa_i_31 : fa_63 port map( a => a(31), b => b(31), ci => carry_s_30_port, co 
                           => c, s => s(31));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity rca_signed_NBIT32_2 is

   port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : out
         std_logic_vector (31 downto 0));

end rca_signed_NBIT32_2;

architecture SYN_Structural of rca_signed_NBIT32_2 is

   component fa_32
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_33
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_34
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_35
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_36
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_37
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_38
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_39
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_40
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_41
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_42
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_43
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_44
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_45
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_46
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_47
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_48
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_49
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_50
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_51
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_52
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_53
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_54
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_55
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_56
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_57
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_58
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_59
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_60
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_61
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_62
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component half_adder_2
      port( a, b : in std_logic;  co, s : out std_logic);
   end component;
   
   signal carry_s_30_port, carry_s_29_port, carry_s_28_port, carry_s_27_port, 
      carry_s_26_port, carry_s_25_port, carry_s_24_port, carry_s_23_port, 
      carry_s_22_port, carry_s_21_port, carry_s_20_port, carry_s_19_port, 
      carry_s_18_port, carry_s_17_port, carry_s_16_port, carry_s_15_port, 
      carry_s_14_port, carry_s_13_port, carry_s_12_port, carry_s_11_port, 
      carry_s_10_port, carry_s_9_port, carry_s_8_port, carry_s_7_port, 
      carry_s_6_port, carry_s_5_port, carry_s_4_port, carry_s_3_port, 
      carry_s_2_port, carry_s_1_port, carry_s_0_port : std_logic;

begin
   
   ha : half_adder_2 port map( a => a(0), b => b(0), co => carry_s_0_port, s =>
                           s(0));
   fa_i_1 : fa_62 port map( a => a(1), b => b(1), ci => carry_s_0_port, co => 
                           carry_s_1_port, s => s(1));
   fa_i_2 : fa_61 port map( a => a(2), b => b(2), ci => carry_s_1_port, co => 
                           carry_s_2_port, s => s(2));
   fa_i_3 : fa_60 port map( a => a(3), b => b(3), ci => carry_s_2_port, co => 
                           carry_s_3_port, s => s(3));
   fa_i_4 : fa_59 port map( a => a(4), b => b(4), ci => carry_s_3_port, co => 
                           carry_s_4_port, s => s(4));
   fa_i_5 : fa_58 port map( a => a(5), b => b(5), ci => carry_s_4_port, co => 
                           carry_s_5_port, s => s(5));
   fa_i_6 : fa_57 port map( a => a(6), b => b(6), ci => carry_s_5_port, co => 
                           carry_s_6_port, s => s(6));
   fa_i_7 : fa_56 port map( a => a(7), b => b(7), ci => carry_s_6_port, co => 
                           carry_s_7_port, s => s(7));
   fa_i_8 : fa_55 port map( a => a(8), b => b(8), ci => carry_s_7_port, co => 
                           carry_s_8_port, s => s(8));
   fa_i_9 : fa_54 port map( a => a(9), b => b(9), ci => carry_s_8_port, co => 
                           carry_s_9_port, s => s(9));
   fa_i_10 : fa_53 port map( a => a(10), b => b(10), ci => carry_s_9_port, co 
                           => carry_s_10_port, s => s(10));
   fa_i_11 : fa_52 port map( a => a(11), b => b(11), ci => carry_s_10_port, co 
                           => carry_s_11_port, s => s(11));
   fa_i_12 : fa_51 port map( a => a(12), b => b(12), ci => carry_s_11_port, co 
                           => carry_s_12_port, s => s(12));
   fa_i_13 : fa_50 port map( a => a(13), b => b(13), ci => carry_s_12_port, co 
                           => carry_s_13_port, s => s(13));
   fa_i_14 : fa_49 port map( a => a(14), b => b(14), ci => carry_s_13_port, co 
                           => carry_s_14_port, s => s(14));
   fa_i_15 : fa_48 port map( a => a(15), b => b(15), ci => carry_s_14_port, co 
                           => carry_s_15_port, s => s(15));
   fa_i_16 : fa_47 port map( a => a(16), b => b(16), ci => carry_s_15_port, co 
                           => carry_s_16_port, s => s(16));
   fa_i_17 : fa_46 port map( a => a(17), b => b(17), ci => carry_s_16_port, co 
                           => carry_s_17_port, s => s(17));
   fa_i_18 : fa_45 port map( a => a(18), b => b(18), ci => carry_s_17_port, co 
                           => carry_s_18_port, s => s(18));
   fa_i_19 : fa_44 port map( a => a(19), b => b(19), ci => carry_s_18_port, co 
                           => carry_s_19_port, s => s(19));
   fa_i_20 : fa_43 port map( a => a(20), b => b(20), ci => carry_s_19_port, co 
                           => carry_s_20_port, s => s(20));
   fa_i_21 : fa_42 port map( a => a(21), b => b(21), ci => carry_s_20_port, co 
                           => carry_s_21_port, s => s(21));
   fa_i_22 : fa_41 port map( a => a(22), b => b(22), ci => carry_s_21_port, co 
                           => carry_s_22_port, s => s(22));
   fa_i_23 : fa_40 port map( a => a(23), b => b(23), ci => carry_s_22_port, co 
                           => carry_s_23_port, s => s(23));
   fa_i_24 : fa_39 port map( a => a(24), b => b(24), ci => carry_s_23_port, co 
                           => carry_s_24_port, s => s(24));
   fa_i_25 : fa_38 port map( a => a(25), b => b(25), ci => carry_s_24_port, co 
                           => carry_s_25_port, s => s(25));
   fa_i_26 : fa_37 port map( a => a(26), b => b(26), ci => carry_s_25_port, co 
                           => carry_s_26_port, s => s(26));
   fa_i_27 : fa_36 port map( a => a(27), b => b(27), ci => carry_s_26_port, co 
                           => carry_s_27_port, s => s(27));
   fa_i_28 : fa_35 port map( a => a(28), b => b(28), ci => carry_s_27_port, co 
                           => carry_s_28_port, s => s(28));
   fa_i_29 : fa_34 port map( a => a(29), b => b(29), ci => carry_s_28_port, co 
                           => carry_s_29_port, s => s(29));
   fa_i_30 : fa_33 port map( a => a(30), b => b(30), ci => carry_s_29_port, co 
                           => carry_s_30_port, s => s(30));
   fa_i_31 : fa_32 port map( a => a(31), b => b(31), ci => carry_s_30_port, co 
                           => c, s => s(31));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity rca_signed_NBIT32_1 is

   port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : out
         std_logic_vector (31 downto 0));

end rca_signed_NBIT32_1;

architecture SYN_Structural of rca_signed_NBIT32_1 is

   component fa_1
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_2
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_3
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_4
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_5
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_6
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_7
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_8
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_9
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_10
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_11
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_12
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_13
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_14
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_15
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_16
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_17
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_18
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_19
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_20
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_21
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_22
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_23
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_24
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_25
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_26
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_27
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_28
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_29
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_30
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_31
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component half_adder_1
      port( a, b : in std_logic;  co, s : out std_logic);
   end component;
   
   signal carry_s_30_port, carry_s_29_port, carry_s_28_port, carry_s_27_port, 
      carry_s_26_port, carry_s_25_port, carry_s_24_port, carry_s_23_port, 
      carry_s_22_port, carry_s_21_port, carry_s_20_port, carry_s_19_port, 
      carry_s_18_port, carry_s_17_port, carry_s_16_port, carry_s_15_port, 
      carry_s_14_port, carry_s_13_port, carry_s_12_port, carry_s_11_port, 
      carry_s_10_port, carry_s_9_port, carry_s_8_port, carry_s_7_port, 
      carry_s_6_port, carry_s_5_port, carry_s_4_port, carry_s_3_port, 
      carry_s_2_port, carry_s_1_port, carry_s_0_port : std_logic;

begin
   
   ha : half_adder_1 port map( a => a(0), b => b(0), co => carry_s_0_port, s =>
                           s(0));
   fa_i_1 : fa_31 port map( a => a(1), b => b(1), ci => carry_s_0_port, co => 
                           carry_s_1_port, s => s(1));
   fa_i_2 : fa_30 port map( a => a(2), b => b(2), ci => carry_s_1_port, co => 
                           carry_s_2_port, s => s(2));
   fa_i_3 : fa_29 port map( a => a(3), b => b(3), ci => carry_s_2_port, co => 
                           carry_s_3_port, s => s(3));
   fa_i_4 : fa_28 port map( a => a(4), b => b(4), ci => carry_s_3_port, co => 
                           carry_s_4_port, s => s(4));
   fa_i_5 : fa_27 port map( a => a(5), b => b(5), ci => carry_s_4_port, co => 
                           carry_s_5_port, s => s(5));
   fa_i_6 : fa_26 port map( a => a(6), b => b(6), ci => carry_s_5_port, co => 
                           carry_s_6_port, s => s(6));
   fa_i_7 : fa_25 port map( a => a(7), b => b(7), ci => carry_s_6_port, co => 
                           carry_s_7_port, s => s(7));
   fa_i_8 : fa_24 port map( a => a(8), b => b(8), ci => carry_s_7_port, co => 
                           carry_s_8_port, s => s(8));
   fa_i_9 : fa_23 port map( a => a(9), b => b(9), ci => carry_s_8_port, co => 
                           carry_s_9_port, s => s(9));
   fa_i_10 : fa_22 port map( a => a(10), b => b(10), ci => carry_s_9_port, co 
                           => carry_s_10_port, s => s(10));
   fa_i_11 : fa_21 port map( a => a(11), b => b(11), ci => carry_s_10_port, co 
                           => carry_s_11_port, s => s(11));
   fa_i_12 : fa_20 port map( a => a(12), b => b(12), ci => carry_s_11_port, co 
                           => carry_s_12_port, s => s(12));
   fa_i_13 : fa_19 port map( a => a(13), b => b(13), ci => carry_s_12_port, co 
                           => carry_s_13_port, s => s(13));
   fa_i_14 : fa_18 port map( a => a(14), b => b(14), ci => carry_s_13_port, co 
                           => carry_s_14_port, s => s(14));
   fa_i_15 : fa_17 port map( a => a(15), b => b(15), ci => carry_s_14_port, co 
                           => carry_s_15_port, s => s(15));
   fa_i_16 : fa_16 port map( a => a(16), b => b(16), ci => carry_s_15_port, co 
                           => carry_s_16_port, s => s(16));
   fa_i_17 : fa_15 port map( a => a(17), b => b(17), ci => carry_s_16_port, co 
                           => carry_s_17_port, s => s(17));
   fa_i_18 : fa_14 port map( a => a(18), b => b(18), ci => carry_s_17_port, co 
                           => carry_s_18_port, s => s(18));
   fa_i_19 : fa_13 port map( a => a(19), b => b(19), ci => carry_s_18_port, co 
                           => carry_s_19_port, s => s(19));
   fa_i_20 : fa_12 port map( a => a(20), b => b(20), ci => carry_s_19_port, co 
                           => carry_s_20_port, s => s(20));
   fa_i_21 : fa_11 port map( a => a(21), b => b(21), ci => carry_s_20_port, co 
                           => carry_s_21_port, s => s(21));
   fa_i_22 : fa_10 port map( a => a(22), b => b(22), ci => carry_s_21_port, co 
                           => carry_s_22_port, s => s(22));
   fa_i_23 : fa_9 port map( a => a(23), b => b(23), ci => carry_s_22_port, co 
                           => carry_s_23_port, s => s(23));
   fa_i_24 : fa_8 port map( a => a(24), b => b(24), ci => carry_s_23_port, co 
                           => carry_s_24_port, s => s(24));
   fa_i_25 : fa_7 port map( a => a(25), b => b(25), ci => carry_s_24_port, co 
                           => carry_s_25_port, s => s(25));
   fa_i_26 : fa_6 port map( a => a(26), b => b(26), ci => carry_s_25_port, co 
                           => carry_s_26_port, s => s(26));
   fa_i_27 : fa_5 port map( a => a(27), b => b(27), ci => carry_s_26_port, co 
                           => carry_s_27_port, s => s(27));
   fa_i_28 : fa_4 port map( a => a(28), b => b(28), ci => carry_s_27_port, co 
                           => carry_s_28_port, s => s(28));
   fa_i_29 : fa_3 port map( a => a(29), b => b(29), ci => carry_s_28_port, co 
                           => carry_s_29_port, s => s(29));
   fa_i_30 : fa_2 port map( a => a(30), b => b(30), ci => carry_s_29_port, co 
                           => carry_s_30_port, s => s(30));
   fa_i_31 : fa_1 port map( a => a(31), b => b(31), ci => carry_s_30_port, co 
                           => c, s => s(31));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_7 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_7;

architecture SYN_behavioral of vp_NBIT32_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U3 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U4 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_6 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_6;

architecture SYN_behavioral of vp_NBIT32_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U3 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U4 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_5 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_5;

architecture SYN_behavioral of vp_NBIT32_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U3 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U4 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_4 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_4;

architecture SYN_behavioral of vp_NBIT32_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U3 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U4 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_3 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_3;

architecture SYN_behavioral of vp_NBIT32_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U3 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U4 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_2 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_2;

architecture SYN_behavioral of vp_NBIT32_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U3 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U4 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_1 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_1;

architecture SYN_behavioral of vp_NBIT32_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U3 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U4 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_7 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_7;

architecture SYN_specification of carry_select_adder_n_bit4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_13
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_14
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_14 port map( operand_1(3) => operand_1(3),
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_13 port map( operand_1(3) => operand_1(3),
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_6 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_6;

architecture SYN_specification of carry_select_adder_n_bit4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_11
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_12
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_12 port map( operand_1(3) => operand_1(3),
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_11 port map( operand_1(3) => operand_1(3),
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_5 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_5;

architecture SYN_specification of carry_select_adder_n_bit4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_9
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_10
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_10 port map( operand_1(3) => operand_1(3),
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_9 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_4 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_4;

architecture SYN_specification of carry_select_adder_n_bit4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_7
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_8
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_8 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_7 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_3 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_3;

architecture SYN_specification of carry_select_adder_n_bit4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_5
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_6
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_6 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_5 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_2 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_2;

architecture SYN_specification of carry_select_adder_n_bit4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_3
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_4
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_4 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_3 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_1 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_1;

architecture SYN_specification of carry_select_adder_n_bit4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_1
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_2
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_2 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_1 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity mux31_N32_1 is

   port( a, b, c : in std_logic_vector (31 downto 0);  sel : in 
         std_logic_vector (1 downto 0);  y : out std_logic_vector (31 downto 0)
         );

end mux31_N32_1;

architecture SYN_Behavioral of mux31_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N37, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15
      , n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35, n36, n37_port, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70 : 
      std_logic;

begin
   
   y_reg_31_inst : DLH_X1 port map( G => N37, D => n70, Q => y(31));
   y_reg_30_inst : DLH_X1 port map( G => N37, D => n69, Q => y(30));
   y_reg_29_inst : DLH_X1 port map( G => N37, D => n68, Q => y(29));
   y_reg_28_inst : DLH_X1 port map( G => N37, D => n67, Q => y(28));
   y_reg_27_inst : DLH_X1 port map( G => N37, D => n66, Q => y(27));
   y_reg_26_inst : DLH_X1 port map( G => N37, D => n65, Q => y(26));
   y_reg_25_inst : DLH_X1 port map( G => N37, D => n64, Q => y(25));
   y_reg_24_inst : DLH_X1 port map( G => N37, D => n63, Q => y(24));
   y_reg_23_inst : DLH_X1 port map( G => N37, D => n62, Q => y(23));
   y_reg_22_inst : DLH_X1 port map( G => N37, D => n61, Q => y(22));
   y_reg_21_inst : DLH_X1 port map( G => N37, D => n60, Q => y(21));
   y_reg_20_inst : DLH_X1 port map( G => N37, D => n59, Q => y(20));
   y_reg_19_inst : DLH_X1 port map( G => N37, D => n58, Q => y(19));
   y_reg_18_inst : DLH_X1 port map( G => N37, D => n57, Q => y(18));
   y_reg_17_inst : DLH_X1 port map( G => N37, D => n56, Q => y(17));
   y_reg_16_inst : DLH_X1 port map( G => N37, D => n55, Q => y(16));
   y_reg_15_inst : DLH_X1 port map( G => N37, D => n54, Q => y(15));
   y_reg_14_inst : DLH_X1 port map( G => N37, D => n53, Q => y(14));
   y_reg_13_inst : DLH_X1 port map( G => N37, D => n52, Q => y(13));
   y_reg_12_inst : DLH_X1 port map( G => N37, D => n51, Q => y(12));
   y_reg_11_inst : DLH_X1 port map( G => N37, D => n50, Q => y(11));
   y_reg_10_inst : DLH_X1 port map( G => N37, D => n49, Q => y(10));
   y_reg_9_inst : DLH_X1 port map( G => N37, D => n48, Q => y(9));
   y_reg_8_inst : DLH_X1 port map( G => N37, D => n47, Q => y(8));
   y_reg_7_inst : DLH_X1 port map( G => N37, D => n46, Q => y(7));
   y_reg_6_inst : DLH_X1 port map( G => N37, D => n45, Q => y(6));
   y_reg_5_inst : DLH_X1 port map( G => N37, D => n44, Q => y(5));
   y_reg_4_inst : DLH_X1 port map( G => N37, D => n43, Q => y(4));
   y_reg_3_inst : DLH_X1 port map( G => N37, D => n42, Q => y(3));
   y_reg_2_inst : DLH_X1 port map( G => N37, D => n41, Q => y(2));
   y_reg_1_inst : DLH_X1 port map( G => N37, D => n40, Q => y(1));
   y_reg_0_inst : DLH_X1 port map( G => N37, D => n39, Q => y(0));
   U3 : OR2_X1 port map( A1 => n3, A2 => n6, ZN => n1);
   U4 : OR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n2);
   U5 : INV_X2 port map( A => n2, ZN => n3);
   U6 : INV_X2 port map( A => n1, ZN => n4);
   U7 : NOR2_X4 port map( A1 => n38, A2 => sel(1), ZN => n6);
   U8 : INV_X1 port map( A => n5, ZN => n39);
   U9 : AOI222_X1 port map( A1 => b(0), A2 => n6, B1 => c(0), B2 => n4, C1 => 
                           a(0), C2 => n3, ZN => n5);
   U10 : INV_X1 port map( A => n7, ZN => n40);
   U11 : AOI222_X1 port map( A1 => b(1), A2 => n6, B1 => c(1), B2 => n4, C1 => 
                           a(1), C2 => n3, ZN => n7);
   U12 : INV_X1 port map( A => n8, ZN => n41);
   U13 : AOI222_X1 port map( A1 => b(2), A2 => n6, B1 => c(2), B2 => n4, C1 => 
                           a(2), C2 => n3, ZN => n8);
   U14 : INV_X1 port map( A => n9, ZN => n42);
   U15 : AOI222_X1 port map( A1 => b(3), A2 => n6, B1 => c(3), B2 => n4, C1 => 
                           a(3), C2 => n3, ZN => n9);
   U16 : INV_X1 port map( A => n10, ZN => n43);
   U17 : AOI222_X1 port map( A1 => b(4), A2 => n6, B1 => c(4), B2 => n4, C1 => 
                           a(4), C2 => n3, ZN => n10);
   U18 : INV_X1 port map( A => n11, ZN => n44);
   U19 : AOI222_X1 port map( A1 => b(5), A2 => n6, B1 => c(5), B2 => n4, C1 => 
                           a(5), C2 => n3, ZN => n11);
   U20 : INV_X1 port map( A => n12, ZN => n45);
   U21 : AOI222_X1 port map( A1 => b(6), A2 => n6, B1 => c(6), B2 => n4, C1 => 
                           a(6), C2 => n3, ZN => n12);
   U22 : INV_X1 port map( A => n13, ZN => n46);
   U23 : AOI222_X1 port map( A1 => b(7), A2 => n6, B1 => c(7), B2 => n4, C1 => 
                           a(7), C2 => n3, ZN => n13);
   U24 : INV_X1 port map( A => n14, ZN => n47);
   U25 : AOI222_X1 port map( A1 => b(8), A2 => n6, B1 => c(8), B2 => n4, C1 => 
                           a(8), C2 => n3, ZN => n14);
   U26 : INV_X1 port map( A => n15, ZN => n48);
   U27 : AOI222_X1 port map( A1 => b(9), A2 => n6, B1 => c(9), B2 => n4, C1 => 
                           a(9), C2 => n3, ZN => n15);
   U28 : INV_X1 port map( A => n16, ZN => n49);
   U29 : AOI222_X1 port map( A1 => b(10), A2 => n6, B1 => c(10), B2 => n4, C1 
                           => a(10), C2 => n3, ZN => n16);
   U30 : INV_X1 port map( A => n17, ZN => n50);
   U31 : AOI222_X1 port map( A1 => b(11), A2 => n6, B1 => c(11), B2 => n4, C1 
                           => a(11), C2 => n3, ZN => n17);
   U32 : INV_X1 port map( A => n18, ZN => n51);
   U33 : AOI222_X1 port map( A1 => b(12), A2 => n6, B1 => c(12), B2 => n4, C1 
                           => a(12), C2 => n3, ZN => n18);
   U34 : INV_X1 port map( A => n19, ZN => n52);
   U35 : AOI222_X1 port map( A1 => b(13), A2 => n6, B1 => c(13), B2 => n4, C1 
                           => a(13), C2 => n3, ZN => n19);
   U36 : INV_X1 port map( A => n20, ZN => n53);
   U37 : AOI222_X1 port map( A1 => b(14), A2 => n6, B1 => c(14), B2 => n4, C1 
                           => a(14), C2 => n3, ZN => n20);
   U38 : INV_X1 port map( A => n21, ZN => n54);
   U39 : AOI222_X1 port map( A1 => b(15), A2 => n6, B1 => c(15), B2 => n4, C1 
                           => a(15), C2 => n3, ZN => n21);
   U40 : INV_X1 port map( A => n22, ZN => n55);
   U41 : AOI222_X1 port map( A1 => b(16), A2 => n6, B1 => c(16), B2 => n4, C1 
                           => a(16), C2 => n3, ZN => n22);
   U42 : INV_X1 port map( A => n23, ZN => n56);
   U43 : AOI222_X1 port map( A1 => b(17), A2 => n6, B1 => c(17), B2 => n4, C1 
                           => a(17), C2 => n3, ZN => n23);
   U44 : INV_X1 port map( A => n24, ZN => n57);
   U45 : AOI222_X1 port map( A1 => b(18), A2 => n6, B1 => c(18), B2 => n4, C1 
                           => a(18), C2 => n3, ZN => n24);
   U46 : INV_X1 port map( A => n25, ZN => n58);
   U47 : AOI222_X1 port map( A1 => b(19), A2 => n6, B1 => c(19), B2 => n4, C1 
                           => a(19), C2 => n3, ZN => n25);
   U48 : INV_X1 port map( A => n26, ZN => n59);
   U49 : AOI222_X1 port map( A1 => b(20), A2 => n6, B1 => c(20), B2 => n4, C1 
                           => a(20), C2 => n3, ZN => n26);
   U50 : INV_X1 port map( A => n27, ZN => n60);
   U51 : AOI222_X1 port map( A1 => b(21), A2 => n6, B1 => c(21), B2 => n4, C1 
                           => a(21), C2 => n3, ZN => n27);
   U52 : INV_X1 port map( A => n28, ZN => n61);
   U53 : AOI222_X1 port map( A1 => b(22), A2 => n6, B1 => c(22), B2 => n4, C1 
                           => a(22), C2 => n3, ZN => n28);
   U54 : INV_X1 port map( A => n29, ZN => n62);
   U55 : AOI222_X1 port map( A1 => b(23), A2 => n6, B1 => c(23), B2 => n4, C1 
                           => a(23), C2 => n3, ZN => n29);
   U56 : INV_X1 port map( A => n30, ZN => n63);
   U57 : AOI222_X1 port map( A1 => b(24), A2 => n6, B1 => c(24), B2 => n4, C1 
                           => a(24), C2 => n3, ZN => n30);
   U58 : INV_X1 port map( A => n31, ZN => n64);
   U59 : AOI222_X1 port map( A1 => b(25), A2 => n6, B1 => c(25), B2 => n4, C1 
                           => a(25), C2 => n3, ZN => n31);
   U60 : INV_X1 port map( A => n32, ZN => n65);
   U61 : AOI222_X1 port map( A1 => b(26), A2 => n6, B1 => c(26), B2 => n4, C1 
                           => a(26), C2 => n3, ZN => n32);
   U62 : INV_X1 port map( A => n33, ZN => n66);
   U63 : AOI222_X1 port map( A1 => b(27), A2 => n6, B1 => c(27), B2 => n4, C1 
                           => a(27), C2 => n3, ZN => n33);
   U64 : INV_X1 port map( A => n34, ZN => n67);
   U65 : AOI222_X1 port map( A1 => b(28), A2 => n6, B1 => c(28), B2 => n4, C1 
                           => a(28), C2 => n3, ZN => n34);
   U66 : INV_X1 port map( A => n35, ZN => n68);
   U67 : AOI222_X1 port map( A1 => b(29), A2 => n6, B1 => c(29), B2 => n4, C1 
                           => a(29), C2 => n3, ZN => n35);
   U68 : INV_X1 port map( A => n36, ZN => n69);
   U69 : AOI222_X1 port map( A1 => b(30), A2 => n6, B1 => c(30), B2 => n4, C1 
                           => a(30), C2 => n3, ZN => n36);
   U70 : INV_X1 port map( A => n37_port, ZN => n70);
   U71 : AOI222_X1 port map( A1 => b(31), A2 => n6, B1 => c(31), B2 => n4, C1 
                           => a(31), C2 => n3, ZN => n37_port);
   U72 : NAND2_X1 port map( A1 => n4, A2 => sel(0), ZN => N37);
   U73 : INV_X1 port map( A => sel(0), ZN => n38);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N5_1 is

   port( a, b : in std_logic_vector (4 downto 0);  sel : in std_logic;  y : out
         std_logic_vector (4 downto 0));

end MUX21_N5_1;

architecture SYN_beh of MUX21_N5_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));
   U2 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U3 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U4 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U5 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N32_6 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end MUX21_N32_6;

architecture SYN_beh of MUX21_N32_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U2 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U3 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U4 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U5 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U6 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U7 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U8 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U9 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U10 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U11 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U12 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U13 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U14 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U15 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U16 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U17 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U18 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U19 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U20 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U21 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U22 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U23 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U24 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U25 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U26 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U27 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U28 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U29 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U30 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U31 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U32 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N32_5 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end MUX21_N32_5;

architecture SYN_beh of MUX21_N32_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U2 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U3 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U4 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U5 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U6 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U7 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U8 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U9 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U10 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U11 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U12 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U13 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U14 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U15 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U16 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U17 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U18 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U19 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U20 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U21 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U22 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U23 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U24 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U25 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U26 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U27 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U28 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U29 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U30 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U31 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U32 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N32_4 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end MUX21_N32_4;

architecture SYN_beh of MUX21_N32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U2 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U3 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U4 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U5 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U6 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U7 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U8 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U9 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U10 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U11 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U12 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U13 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U14 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U15 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U16 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U17 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U18 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U19 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U20 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U21 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U22 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U23 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U24 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U25 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U26 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U27 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U28 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U29 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U30 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U31 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U32 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N32_3 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end MUX21_N32_3;

architecture SYN_beh of MUX21_N32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U2 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U3 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U4 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U5 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U6 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U7 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U8 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U9 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U10 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U11 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U12 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U13 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U14 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U15 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U16 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U17 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U18 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U19 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U20 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U21 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U22 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U23 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U24 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U25 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U26 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U27 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U28 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U29 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U30 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U31 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U32 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N32_2 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end MUX21_N32_2;

architecture SYN_beh of MUX21_N32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));
   U2 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U3 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U4 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U5 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U6 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U7 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U8 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U9 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U10 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U11 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U12 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U13 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U14 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U15 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U16 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U17 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U18 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U19 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U20 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U21 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U22 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U23 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U24 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U25 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U26 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U27 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U28 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U29 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U30 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U31 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U32 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N32_1 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end MUX21_N32_1;

architecture SYN_beh of MUX21_N32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U2 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U3 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U4 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U5 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U6 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U7 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U8 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U9 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U10 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U11 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U12 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U13 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U14 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U15 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U16 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U17 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U18 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U19 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U20 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U21 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U22 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U23 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U24 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U25 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U26 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U27 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U28 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U29 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U30 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U31 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U32 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity or2_0 is

   port( a, b : in std_logic;  o : out std_logic);

end or2_0;

architecture SYN_Behavioral of or2_0 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => a, A2 => b, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity xor2_0 is

   port( a, b : in std_logic;  o : out std_logic);

end xor2_0;

architecture SYN_Behavioral of xor2_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity and2_0 is

   port( a, b : in std_logic;  o : out std_logic);

end and2_0;

architecture SYN_Behavioral of and2_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => o);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity full_adder_0 is

   port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : out 
         std_logic);

end full_adder_0;

architecture SYN_full_adder_arc of full_adder_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => carry_in, B => n1, Z => sum);
   U2 : INV_X1 port map( A => n2, ZN => carry_out);
   U3 : AOI22_X1 port map( A1 => operand_2, A2 => operand_1, B1 => n1, B2 => 
                           carry_in, ZN => n2);
   U4 : XOR2_X1 port map( A => operand_1, B => operand_2, Z => n1);

end SYN_full_adder_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fa_0 is

   port( a, b, ci : in std_logic;  co, s : out std_logic);

end fa_0;

architecture SYN_Structural of fa_0 is

   component or2_0
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_439
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_440
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_439
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component xor2_440
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   signal s1, s2, s3 : std_logic;

begin
   
   xor_1 : xor2_440 port map( a => a, b => b, o => s1);
   xor_2 : xor2_439 port map( a => s1, b => ci, o => s);
   and_1 : and2_440 port map( a => a, b => b, o => s2);
   and_2 : and2_439 port map( a => s1, b => ci, o => s3);
   or_1 : or2_0 port map( a => s2, b => s3, o => co);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity half_adder_0 is

   port( a, b : in std_logic;  co, s : out std_logic);

end half_adder_0;

architecture SYN_Structural of half_adder_0 is

   component xor2_0
      port( a, b : in std_logic;  o : out std_logic);
   end component;
   
   component and2_0
      port( a, b : in std_logic;  o : out std_logic);
   end component;

begin
   
   carry : and2_0 port map( a => a, b => b, o => co);
   sum : xor2_0 port map( a => a, b => b, o => s);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ripple_carry_adder_n_bit4_0 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end ripple_carry_adder_n_bit4_0;

architecture SYN_rca_arc of ripple_carry_adder_n_bit4_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component full_adder_61
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_62
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_63
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   component full_adder_0
      port( operand_1, operand_2, carry_in : in std_logic;  sum, carry_out : 
            out std_logic);
   end component;
   
   signal carry_out_port, cin_3_port, cin_2_port, cin_1_port : std_logic;

begin
   carry_out <= carry_out_port;
   
   f_adder_0 : full_adder_0 port map( operand_1 => operand_1(0), operand_2 => 
                           operand_2(0), carry_in => carry_in, sum => sum(0), 
                           carry_out => cin_1_port);
   f_adder_1 : full_adder_63 port map( operand_1 => operand_1(1), operand_2 => 
                           operand_2(1), carry_in => cin_1_port, sum => sum(1),
                           carry_out => cin_2_port);
   f_adder_2 : full_adder_62 port map( operand_1 => operand_1(2), operand_2 => 
                           operand_2(2), carry_in => cin_2_port, sum => sum(2),
                           carry_out => cin_3_port);
   f_adder_3 : full_adder_61 port map( operand_1 => operand_1(3), operand_2 => 
                           operand_2(3), carry_in => cin_3_port, sum => sum(3),
                           carry_out => carry_out_port);
   U1 : XOR2_X1 port map( A => cin_3_port, B => carry_out_port, Z => overflow);

end SYN_rca_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_0 is

   port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);

end g_block_0;

architecture SYN_specification of g_block_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_block_0 is

   port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);

end pg_block_0;

architecture SYN_specification of pg_block_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk1j, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pk1j, A2 => Pik, ZN => Pij);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity g_block_carry is

   port( Gik, Pik, Gk1j, Pk1j, carry_in : in std_logic;  Gij : out std_logic);

end g_block_carry;

architecture SYN_specification of g_block_carry is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => Gij);
   U2 : INV_X1 port map( A => Gik, ZN => n3);
   U3 : INV_X1 port map( A => Pik, ZN => n2);
   U4 : AOI21_X1 port map( B1 => carry_in, B2 => Pk1j, A => Gk1j, ZN => n1);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity pg_network_n_bit32 is

   port( operand_1, operand_2 : in std_logic_vector (32 downto 1);  p, g : out 
         std_logic_vector (32 downto 1));

end pg_network_n_bit32;

architecture SYN_specification of pg_network_n_bit32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => operand_2(9), B => operand_1(9), Z => p(9));
   U2 : XOR2_X1 port map( A => operand_2(8), B => operand_1(8), Z => p(8));
   U3 : XOR2_X1 port map( A => operand_2(7), B => operand_1(7), Z => p(7));
   U4 : XOR2_X1 port map( A => operand_2(6), B => operand_1(6), Z => p(6));
   U5 : XOR2_X1 port map( A => operand_2(5), B => operand_1(5), Z => p(5));
   U6 : XOR2_X1 port map( A => operand_2(4), B => operand_1(4), Z => p(4));
   U7 : XOR2_X1 port map( A => operand_2(3), B => operand_1(3), Z => p(3));
   U8 : XOR2_X1 port map( A => operand_2(32), B => operand_1(32), Z => p(32));
   U9 : XOR2_X1 port map( A => operand_2(31), B => operand_1(31), Z => p(31));
   U10 : XOR2_X1 port map( A => operand_2(30), B => operand_1(30), Z => p(30));
   U11 : XOR2_X1 port map( A => operand_2(2), B => operand_1(2), Z => p(2));
   U12 : XOR2_X1 port map( A => operand_2(29), B => operand_1(29), Z => p(29));
   U13 : XOR2_X1 port map( A => operand_2(28), B => operand_1(28), Z => p(28));
   U14 : XOR2_X1 port map( A => operand_2(27), B => operand_1(27), Z => p(27));
   U15 : XOR2_X1 port map( A => operand_2(26), B => operand_1(26), Z => p(26));
   U16 : XOR2_X1 port map( A => operand_2(25), B => operand_1(25), Z => p(25));
   U17 : XOR2_X1 port map( A => operand_2(24), B => operand_1(24), Z => p(24));
   U18 : XOR2_X1 port map( A => operand_2(23), B => operand_1(23), Z => p(23));
   U19 : XOR2_X1 port map( A => operand_2(22), B => operand_1(22), Z => p(22));
   U20 : XOR2_X1 port map( A => operand_2(21), B => operand_1(21), Z => p(21));
   U21 : XOR2_X1 port map( A => operand_2(20), B => operand_1(20), Z => p(20));
   U22 : XOR2_X1 port map( A => operand_2(1), B => operand_1(1), Z => p(1));
   U23 : XOR2_X1 port map( A => operand_2(19), B => operand_1(19), Z => p(19));
   U24 : XOR2_X1 port map( A => operand_2(18), B => operand_1(18), Z => p(18));
   U25 : XOR2_X1 port map( A => operand_2(17), B => operand_1(17), Z => p(17));
   U26 : XOR2_X1 port map( A => operand_2(16), B => operand_1(16), Z => p(16));
   U27 : XOR2_X1 port map( A => operand_2(15), B => operand_1(15), Z => p(15));
   U28 : XOR2_X1 port map( A => operand_2(14), B => operand_1(14), Z => p(14));
   U29 : XOR2_X1 port map( A => operand_2(13), B => operand_1(13), Z => p(13));
   U30 : XOR2_X1 port map( A => operand_2(12), B => operand_1(12), Z => p(12));
   U31 : XOR2_X1 port map( A => operand_2(11), B => operand_1(11), Z => p(11));
   U32 : XOR2_X1 port map( A => operand_2(10), B => operand_1(10), Z => p(10));
   U33 : AND2_X1 port map( A1 => operand_2(9), A2 => operand_1(9), ZN => g(9));
   U34 : AND2_X1 port map( A1 => operand_2(8), A2 => operand_1(8), ZN => g(8));
   U35 : AND2_X1 port map( A1 => operand_2(7), A2 => operand_1(7), ZN => g(7));
   U36 : AND2_X1 port map( A1 => operand_2(6), A2 => operand_1(6), ZN => g(6));
   U37 : AND2_X1 port map( A1 => operand_2(5), A2 => operand_1(5), ZN => g(5));
   U38 : AND2_X1 port map( A1 => operand_2(4), A2 => operand_1(4), ZN => g(4));
   U39 : AND2_X1 port map( A1 => operand_2(3), A2 => operand_1(3), ZN => g(3));
   U40 : AND2_X1 port map( A1 => operand_2(32), A2 => operand_1(32), ZN => 
                           g(32));
   U41 : AND2_X1 port map( A1 => operand_2(31), A2 => operand_1(31), ZN => 
                           g(31));
   U42 : AND2_X1 port map( A1 => operand_2(30), A2 => operand_1(30), ZN => 
                           g(30));
   U43 : AND2_X1 port map( A1 => operand_2(2), A2 => operand_1(2), ZN => g(2));
   U44 : AND2_X1 port map( A1 => operand_2(29), A2 => operand_1(29), ZN => 
                           g(29));
   U45 : AND2_X1 port map( A1 => operand_2(28), A2 => operand_1(28), ZN => 
                           g(28));
   U46 : AND2_X1 port map( A1 => operand_2(27), A2 => operand_1(27), ZN => 
                           g(27));
   U47 : AND2_X1 port map( A1 => operand_2(26), A2 => operand_1(26), ZN => 
                           g(26));
   U48 : AND2_X1 port map( A1 => operand_2(25), A2 => operand_1(25), ZN => 
                           g(25));
   U49 : AND2_X1 port map( A1 => operand_2(24), A2 => operand_1(24), ZN => 
                           g(24));
   U50 : AND2_X1 port map( A1 => operand_2(23), A2 => operand_1(23), ZN => 
                           g(23));
   U51 : AND2_X1 port map( A1 => operand_2(22), A2 => operand_1(22), ZN => 
                           g(22));
   U52 : AND2_X1 port map( A1 => operand_2(21), A2 => operand_1(21), ZN => 
                           g(21));
   U53 : AND2_X1 port map( A1 => operand_2(20), A2 => operand_1(20), ZN => 
                           g(20));
   U54 : AND2_X1 port map( A1 => operand_2(1), A2 => operand_1(1), ZN => g(1));
   U55 : AND2_X1 port map( A1 => operand_2(19), A2 => operand_1(19), ZN => 
                           g(19));
   U56 : AND2_X1 port map( A1 => operand_2(18), A2 => operand_1(18), ZN => 
                           g(18));
   U57 : AND2_X1 port map( A1 => operand_2(17), A2 => operand_1(17), ZN => 
                           g(17));
   U58 : AND2_X1 port map( A1 => operand_2(16), A2 => operand_1(16), ZN => 
                           g(16));
   U59 : AND2_X1 port map( A1 => operand_2(15), A2 => operand_1(15), ZN => 
                           g(15));
   U60 : AND2_X1 port map( A1 => operand_2(14), A2 => operand_1(14), ZN => 
                           g(14));
   U61 : AND2_X1 port map( A1 => operand_2(13), A2 => operand_1(13), ZN => 
                           g(13));
   U62 : AND2_X1 port map( A1 => operand_2(12), A2 => operand_1(12), ZN => 
                           g(12));
   U63 : AND2_X1 port map( A1 => operand_2(11), A2 => operand_1(11), ZN => 
                           g(11));
   U64 : AND2_X1 port map( A1 => operand_2(10), A2 => operand_1(10), ZN => 
                           g(10));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX81_N32 is

   port( a, b, c, d, e, f, g, h : in std_logic_vector (31 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32;

architecture SYN_beh of MUX81_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148 : std_logic;

begin
   
   U1 : OR4_X1 port map( A1 => n9, A2 => n4, A3 => n3, A4 => n145, ZN => n1);
   U2 : INV_X2 port map( A => n1, ZN => n2);
   U3 : OR3_X1 port map( A1 => sel(1), A2 => sel(2), A3 => n146, ZN => n14);
   U4 : INV_X2 port map( A => n14, ZN => n3);
   U5 : OR3_X1 port map( A1 => n147, A2 => sel(0), A3 => n148, ZN => n16);
   U6 : INV_X2 port map( A => n16, ZN => n4);
   U7 : OR3_X1 port map( A1 => sel(0), A2 => sel(2), A3 => n147, ZN => n18);
   U8 : INV_X2 port map( A => n18, ZN => n5);
   U9 : OR3_X1 port map( A1 => n146, A2 => sel(1), A3 => n148, ZN => n17);
   U10 : INV_X2 port map( A => n17, ZN => n6);
   U11 : OR3_X1 port map( A1 => sel(1), A2 => sel(2), A3 => sel(0), ZN => n19);
   U12 : INV_X2 port map( A => n19, ZN => n7);
   U13 : OR3_X1 port map( A1 => n146, A2 => sel(2), A3 => n147, ZN => n20);
   U14 : INV_X2 port map( A => n20, ZN => n8);
   U15 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n148, ZN => n15);
   U16 : INV_X2 port map( A => n15, ZN => n9);
   U17 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => 
                           y(9));
   U18 : AOI22_X1 port map( A1 => h(9), A2 => n2, B1 => b(9), B2 => n3, ZN => 
                           n13);
   U19 : AOI22_X1 port map( A1 => e(9), A2 => n9, B1 => g(9), B2 => n4, ZN => 
                           n12);
   U20 : AOI22_X1 port map( A1 => f(9), A2 => n6, B1 => c(9), B2 => n5, ZN => 
                           n11);
   U21 : AOI22_X1 port map( A1 => a(9), A2 => n7, B1 => d(9), B2 => n8, ZN => 
                           n10);
   U22 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           y(8));
   U23 : AOI22_X1 port map( A1 => h(8), A2 => n2, B1 => b(8), B2 => n3, ZN => 
                           n24);
   U24 : AOI22_X1 port map( A1 => e(8), A2 => n9, B1 => g(8), B2 => n4, ZN => 
                           n23);
   U25 : AOI22_X1 port map( A1 => f(8), A2 => n6, B1 => c(8), B2 => n5, ZN => 
                           n22);
   U26 : AOI22_X1 port map( A1 => a(8), A2 => n7, B1 => d(8), B2 => n8, ZN => 
                           n21);
   U27 : NAND4_X1 port map( A1 => n25, A2 => n26, A3 => n27, A4 => n28, ZN => 
                           y(7));
   U28 : AOI22_X1 port map( A1 => h(7), A2 => n2, B1 => b(7), B2 => n3, ZN => 
                           n28);
   U29 : AOI22_X1 port map( A1 => e(7), A2 => n9, B1 => g(7), B2 => n4, ZN => 
                           n27);
   U30 : AOI22_X1 port map( A1 => f(7), A2 => n6, B1 => c(7), B2 => n5, ZN => 
                           n26);
   U31 : AOI22_X1 port map( A1 => a(7), A2 => n7, B1 => d(7), B2 => n8, ZN => 
                           n25);
   U32 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           y(6));
   U33 : AOI22_X1 port map( A1 => h(6), A2 => n2, B1 => b(6), B2 => n3, ZN => 
                           n32);
   U34 : AOI22_X1 port map( A1 => e(6), A2 => n9, B1 => g(6), B2 => n4, ZN => 
                           n31);
   U35 : AOI22_X1 port map( A1 => f(6), A2 => n6, B1 => c(6), B2 => n5, ZN => 
                           n30);
   U36 : AOI22_X1 port map( A1 => a(6), A2 => n7, B1 => d(6), B2 => n8, ZN => 
                           n29);
   U37 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           y(5));
   U38 : AOI22_X1 port map( A1 => h(5), A2 => n2, B1 => b(5), B2 => n3, ZN => 
                           n36);
   U39 : AOI22_X1 port map( A1 => e(5), A2 => n9, B1 => g(5), B2 => n4, ZN => 
                           n35);
   U40 : AOI22_X1 port map( A1 => f(5), A2 => n6, B1 => c(5), B2 => n5, ZN => 
                           n34);
   U41 : AOI22_X1 port map( A1 => a(5), A2 => n7, B1 => d(5), B2 => n8, ZN => 
                           n33);
   U42 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           y(4));
   U43 : AOI22_X1 port map( A1 => h(4), A2 => n2, B1 => b(4), B2 => n3, ZN => 
                           n40);
   U44 : AOI22_X1 port map( A1 => e(4), A2 => n9, B1 => g(4), B2 => n4, ZN => 
                           n39);
   U45 : AOI22_X1 port map( A1 => f(4), A2 => n6, B1 => c(4), B2 => n5, ZN => 
                           n38);
   U46 : AOI22_X1 port map( A1 => a(4), A2 => n7, B1 => d(4), B2 => n8, ZN => 
                           n37);
   U47 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           y(3));
   U48 : AOI22_X1 port map( A1 => h(3), A2 => n2, B1 => b(3), B2 => n3, ZN => 
                           n44);
   U49 : AOI22_X1 port map( A1 => e(3), A2 => n9, B1 => g(3), B2 => n4, ZN => 
                           n43);
   U50 : AOI22_X1 port map( A1 => f(3), A2 => n6, B1 => c(3), B2 => n5, ZN => 
                           n42);
   U51 : AOI22_X1 port map( A1 => a(3), A2 => n7, B1 => d(3), B2 => n8, ZN => 
                           n41);
   U52 : NAND4_X1 port map( A1 => n45, A2 => n46, A3 => n47, A4 => n48, ZN => 
                           y(31));
   U53 : AOI22_X1 port map( A1 => h(31), A2 => n2, B1 => b(31), B2 => n3, ZN =>
                           n48);
   U54 : AOI22_X1 port map( A1 => e(31), A2 => n9, B1 => g(31), B2 => n4, ZN =>
                           n47);
   U55 : AOI22_X1 port map( A1 => f(31), A2 => n6, B1 => c(31), B2 => n5, ZN =>
                           n46);
   U56 : AOI22_X1 port map( A1 => a(31), A2 => n7, B1 => d(31), B2 => n8, ZN =>
                           n45);
   U57 : NAND4_X1 port map( A1 => n49, A2 => n50, A3 => n51, A4 => n52, ZN => 
                           y(30));
   U58 : AOI22_X1 port map( A1 => h(30), A2 => n2, B1 => b(30), B2 => n3, ZN =>
                           n52);
   U59 : AOI22_X1 port map( A1 => e(30), A2 => n9, B1 => g(30), B2 => n4, ZN =>
                           n51);
   U60 : AOI22_X1 port map( A1 => f(30), A2 => n6, B1 => c(30), B2 => n5, ZN =>
                           n50);
   U61 : AOI22_X1 port map( A1 => a(30), A2 => n7, B1 => d(30), B2 => n8, ZN =>
                           n49);
   U62 : NAND4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           y(2));
   U63 : AOI22_X1 port map( A1 => h(2), A2 => n2, B1 => b(2), B2 => n3, ZN => 
                           n56);
   U64 : AOI22_X1 port map( A1 => e(2), A2 => n9, B1 => g(2), B2 => n4, ZN => 
                           n55);
   U65 : AOI22_X1 port map( A1 => f(2), A2 => n6, B1 => c(2), B2 => n5, ZN => 
                           n54);
   U66 : AOI22_X1 port map( A1 => a(2), A2 => n7, B1 => d(2), B2 => n8, ZN => 
                           n53);
   U67 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           y(29));
   U68 : AOI22_X1 port map( A1 => h(29), A2 => n2, B1 => b(29), B2 => n3, ZN =>
                           n60);
   U69 : AOI22_X1 port map( A1 => e(29), A2 => n9, B1 => g(29), B2 => n4, ZN =>
                           n59);
   U70 : AOI22_X1 port map( A1 => f(29), A2 => n6, B1 => c(29), B2 => n5, ZN =>
                           n58);
   U71 : AOI22_X1 port map( A1 => a(29), A2 => n7, B1 => d(29), B2 => n8, ZN =>
                           n57);
   U72 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           y(28));
   U73 : AOI22_X1 port map( A1 => h(28), A2 => n2, B1 => b(28), B2 => n3, ZN =>
                           n64);
   U74 : AOI22_X1 port map( A1 => e(28), A2 => n9, B1 => g(28), B2 => n4, ZN =>
                           n63);
   U75 : AOI22_X1 port map( A1 => f(28), A2 => n6, B1 => c(28), B2 => n5, ZN =>
                           n62);
   U76 : AOI22_X1 port map( A1 => a(28), A2 => n7, B1 => d(28), B2 => n8, ZN =>
                           n61);
   U77 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           y(27));
   U78 : AOI22_X1 port map( A1 => h(27), A2 => n2, B1 => b(27), B2 => n3, ZN =>
                           n68);
   U79 : AOI22_X1 port map( A1 => e(27), A2 => n9, B1 => g(27), B2 => n4, ZN =>
                           n67);
   U80 : AOI22_X1 port map( A1 => f(27), A2 => n6, B1 => c(27), B2 => n5, ZN =>
                           n66);
   U81 : AOI22_X1 port map( A1 => a(27), A2 => n7, B1 => d(27), B2 => n8, ZN =>
                           n65);
   U82 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           y(26));
   U83 : AOI22_X1 port map( A1 => h(26), A2 => n2, B1 => b(26), B2 => n3, ZN =>
                           n72);
   U84 : AOI22_X1 port map( A1 => e(26), A2 => n9, B1 => g(26), B2 => n4, ZN =>
                           n71);
   U85 : AOI22_X1 port map( A1 => f(26), A2 => n6, B1 => c(26), B2 => n5, ZN =>
                           n70);
   U86 : AOI22_X1 port map( A1 => a(26), A2 => n7, B1 => d(26), B2 => n8, ZN =>
                           n69);
   U87 : NAND4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           y(25));
   U88 : AOI22_X1 port map( A1 => h(25), A2 => n2, B1 => b(25), B2 => n3, ZN =>
                           n76);
   U89 : AOI22_X1 port map( A1 => e(25), A2 => n9, B1 => g(25), B2 => n4, ZN =>
                           n75);
   U90 : AOI22_X1 port map( A1 => f(25), A2 => n6, B1 => c(25), B2 => n5, ZN =>
                           n74);
   U91 : AOI22_X1 port map( A1 => a(25), A2 => n7, B1 => d(25), B2 => n8, ZN =>
                           n73);
   U92 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           y(24));
   U93 : AOI22_X1 port map( A1 => h(24), A2 => n2, B1 => b(24), B2 => n3, ZN =>
                           n80);
   U94 : AOI22_X1 port map( A1 => e(24), A2 => n9, B1 => g(24), B2 => n4, ZN =>
                           n79);
   U95 : AOI22_X1 port map( A1 => f(24), A2 => n6, B1 => c(24), B2 => n5, ZN =>
                           n78);
   U96 : AOI22_X1 port map( A1 => a(24), A2 => n7, B1 => d(24), B2 => n8, ZN =>
                           n77);
   U97 : NAND4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           y(23));
   U98 : AOI22_X1 port map( A1 => h(23), A2 => n2, B1 => b(23), B2 => n3, ZN =>
                           n84);
   U99 : AOI22_X1 port map( A1 => e(23), A2 => n9, B1 => g(23), B2 => n4, ZN =>
                           n83);
   U100 : AOI22_X1 port map( A1 => f(23), A2 => n6, B1 => c(23), B2 => n5, ZN 
                           => n82);
   U101 : AOI22_X1 port map( A1 => a(23), A2 => n7, B1 => d(23), B2 => n8, ZN 
                           => n81);
   U102 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           y(22));
   U103 : AOI22_X1 port map( A1 => h(22), A2 => n2, B1 => b(22), B2 => n3, ZN 
                           => n88);
   U104 : AOI22_X1 port map( A1 => e(22), A2 => n9, B1 => g(22), B2 => n4, ZN 
                           => n87);
   U105 : AOI22_X1 port map( A1 => f(22), A2 => n6, B1 => c(22), B2 => n5, ZN 
                           => n86);
   U106 : AOI22_X1 port map( A1 => a(22), A2 => n7, B1 => d(22), B2 => n8, ZN 
                           => n85);
   U107 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           y(21));
   U108 : AOI22_X1 port map( A1 => h(21), A2 => n2, B1 => b(21), B2 => n3, ZN 
                           => n92);
   U109 : AOI22_X1 port map( A1 => e(21), A2 => n9, B1 => g(21), B2 => n4, ZN 
                           => n91);
   U110 : AOI22_X1 port map( A1 => f(21), A2 => n6, B1 => c(21), B2 => n5, ZN 
                           => n90);
   U111 : AOI22_X1 port map( A1 => a(21), A2 => n7, B1 => d(21), B2 => n8, ZN 
                           => n89);
   U112 : NAND4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           y(20));
   U113 : AOI22_X1 port map( A1 => h(20), A2 => n2, B1 => b(20), B2 => n3, ZN 
                           => n96);
   U114 : AOI22_X1 port map( A1 => e(20), A2 => n9, B1 => g(20), B2 => n4, ZN 
                           => n95);
   U115 : AOI22_X1 port map( A1 => f(20), A2 => n6, B1 => c(20), B2 => n5, ZN 
                           => n94);
   U116 : AOI22_X1 port map( A1 => a(20), A2 => n7, B1 => d(20), B2 => n8, ZN 
                           => n93);
   U117 : NAND4_X1 port map( A1 => n97, A2 => n98, A3 => n99, A4 => n100, ZN =>
                           y(1));
   U118 : AOI22_X1 port map( A1 => h(1), A2 => n2, B1 => b(1), B2 => n3, ZN => 
                           n100);
   U119 : AOI22_X1 port map( A1 => e(1), A2 => n9, B1 => g(1), B2 => n4, ZN => 
                           n99);
   U120 : AOI22_X1 port map( A1 => f(1), A2 => n6, B1 => c(1), B2 => n5, ZN => 
                           n98);
   U121 : AOI22_X1 port map( A1 => a(1), A2 => n7, B1 => d(1), B2 => n8, ZN => 
                           n97);
   U122 : NAND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN
                           => y(19));
   U123 : AOI22_X1 port map( A1 => h(19), A2 => n2, B1 => b(19), B2 => n3, ZN 
                           => n104);
   U124 : AOI22_X1 port map( A1 => e(19), A2 => n9, B1 => g(19), B2 => n4, ZN 
                           => n103);
   U125 : AOI22_X1 port map( A1 => f(19), A2 => n6, B1 => c(19), B2 => n5, ZN 
                           => n102);
   U126 : AOI22_X1 port map( A1 => a(19), A2 => n7, B1 => d(19), B2 => n8, ZN 
                           => n101);
   U127 : NAND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN
                           => y(18));
   U128 : AOI22_X1 port map( A1 => h(18), A2 => n2, B1 => b(18), B2 => n3, ZN 
                           => n108);
   U129 : AOI22_X1 port map( A1 => e(18), A2 => n9, B1 => g(18), B2 => n4, ZN 
                           => n107);
   U130 : AOI22_X1 port map( A1 => f(18), A2 => n6, B1 => c(18), B2 => n5, ZN 
                           => n106);
   U131 : AOI22_X1 port map( A1 => a(18), A2 => n7, B1 => d(18), B2 => n8, ZN 
                           => n105);
   U132 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => y(17));
   U133 : AOI22_X1 port map( A1 => h(17), A2 => n2, B1 => b(17), B2 => n3, ZN 
                           => n112);
   U134 : AOI22_X1 port map( A1 => e(17), A2 => n9, B1 => g(17), B2 => n4, ZN 
                           => n111);
   U135 : AOI22_X1 port map( A1 => f(17), A2 => n6, B1 => c(17), B2 => n5, ZN 
                           => n110);
   U136 : AOI22_X1 port map( A1 => a(17), A2 => n7, B1 => d(17), B2 => n8, ZN 
                           => n109);
   U137 : NAND4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN
                           => y(16));
   U138 : AOI22_X1 port map( A1 => h(16), A2 => n2, B1 => b(16), B2 => n3, ZN 
                           => n116);
   U139 : AOI22_X1 port map( A1 => e(16), A2 => n9, B1 => g(16), B2 => n4, ZN 
                           => n115);
   U140 : AOI22_X1 port map( A1 => f(16), A2 => n6, B1 => c(16), B2 => n5, ZN 
                           => n114);
   U141 : AOI22_X1 port map( A1 => a(16), A2 => n7, B1 => d(16), B2 => n8, ZN 
                           => n113);
   U142 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN
                           => y(15));
   U143 : AOI22_X1 port map( A1 => h(15), A2 => n2, B1 => b(15), B2 => n3, ZN 
                           => n120);
   U144 : AOI22_X1 port map( A1 => e(15), A2 => n9, B1 => g(15), B2 => n4, ZN 
                           => n119);
   U145 : AOI22_X1 port map( A1 => f(15), A2 => n6, B1 => c(15), B2 => n5, ZN 
                           => n118);
   U146 : AOI22_X1 port map( A1 => a(15), A2 => n7, B1 => d(15), B2 => n8, ZN 
                           => n117);
   U147 : NAND4_X1 port map( A1 => n121, A2 => n122, A3 => n123, A4 => n124, ZN
                           => y(14));
   U148 : AOI22_X1 port map( A1 => h(14), A2 => n2, B1 => b(14), B2 => n3, ZN 
                           => n124);
   U149 : AOI22_X1 port map( A1 => e(14), A2 => n9, B1 => g(14), B2 => n4, ZN 
                           => n123);
   U150 : AOI22_X1 port map( A1 => f(14), A2 => n6, B1 => c(14), B2 => n5, ZN 
                           => n122);
   U151 : AOI22_X1 port map( A1 => a(14), A2 => n7, B1 => d(14), B2 => n8, ZN 
                           => n121);
   U152 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => y(13));
   U153 : AOI22_X1 port map( A1 => h(13), A2 => n2, B1 => b(13), B2 => n3, ZN 
                           => n128);
   U154 : AOI22_X1 port map( A1 => e(13), A2 => n9, B1 => g(13), B2 => n4, ZN 
                           => n127);
   U155 : AOI22_X1 port map( A1 => f(13), A2 => n6, B1 => c(13), B2 => n5, ZN 
                           => n126);
   U156 : AOI22_X1 port map( A1 => a(13), A2 => n7, B1 => d(13), B2 => n8, ZN 
                           => n125);
   U157 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => y(12));
   U158 : AOI22_X1 port map( A1 => h(12), A2 => n2, B1 => b(12), B2 => n3, ZN 
                           => n132);
   U159 : AOI22_X1 port map( A1 => e(12), A2 => n9, B1 => g(12), B2 => n4, ZN 
                           => n131);
   U160 : AOI22_X1 port map( A1 => f(12), A2 => n6, B1 => c(12), B2 => n5, ZN 
                           => n130);
   U161 : AOI22_X1 port map( A1 => a(12), A2 => n7, B1 => d(12), B2 => n8, ZN 
                           => n129);
   U162 : NAND4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN
                           => y(11));
   U163 : AOI22_X1 port map( A1 => h(11), A2 => n2, B1 => b(11), B2 => n3, ZN 
                           => n136);
   U164 : AOI22_X1 port map( A1 => e(11), A2 => n9, B1 => g(11), B2 => n4, ZN 
                           => n135);
   U165 : AOI22_X1 port map( A1 => f(11), A2 => n6, B1 => c(11), B2 => n5, ZN 
                           => n134);
   U166 : AOI22_X1 port map( A1 => a(11), A2 => n7, B1 => d(11), B2 => n8, ZN 
                           => n133);
   U167 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => y(10));
   U168 : AOI22_X1 port map( A1 => h(10), A2 => n2, B1 => b(10), B2 => n3, ZN 
                           => n140);
   U169 : AOI22_X1 port map( A1 => e(10), A2 => n9, B1 => g(10), B2 => n4, ZN 
                           => n139);
   U170 : AOI22_X1 port map( A1 => f(10), A2 => n6, B1 => c(10), B2 => n5, ZN 
                           => n138);
   U171 : AOI22_X1 port map( A1 => a(10), A2 => n7, B1 => d(10), B2 => n8, ZN 
                           => n137);
   U172 : NAND4_X1 port map( A1 => n141, A2 => n142, A3 => n143, A4 => n144, ZN
                           => y(0));
   U173 : AOI22_X1 port map( A1 => h(0), A2 => n2, B1 => b(0), B2 => n3, ZN => 
                           n144);
   U174 : OR4_X1 port map( A1 => n8, A2 => n7, A3 => n5, A4 => n6, ZN => n145);
   U175 : AOI22_X1 port map( A1 => e(0), A2 => n9, B1 => g(0), B2 => n4, ZN => 
                           n143);
   U176 : AOI22_X1 port map( A1 => f(0), A2 => n6, B1 => c(0), B2 => n5, ZN => 
                           n142);
   U177 : INV_X1 port map( A => sel(2), ZN => n148);
   U178 : AOI22_X1 port map( A1 => a(0), A2 => n7, B1 => d(0), B2 => n8, ZN => 
                           n141);
   U179 : INV_X1 port map( A => sel(1), ZN => n147);
   U180 : INV_X1 port map( A => sel(0), ZN => n146);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX41_N40 is

   port( a, b, c, d : in std_logic_vector (39 downto 0);  sel : in 
         std_logic_vector (1 downto 0);  y : out std_logic_vector (39 downto 0)
         );

end MUX41_N40;

architecture SYN_beh of MUX41_N40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86 : std_logic;

begin
   
   U1 : CLKBUF_X2 port map( A => n4, Z => n1);
   U2 : NOR2_X4 port map( A1 => n86, A2 => sel(0), ZN => n7);
   U3 : AND2_X2 port map( A1 => sel(0), A2 => n86, ZN => n5);
   U4 : NOR2_X4 port map( A1 => sel(0), A2 => sel(1), ZN => n6);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => y(9));
   U6 : AOI22_X1 port map( A1 => d(9), A2 => n1, B1 => b(9), B2 => n5, ZN => n3
                           );
   U7 : AOI22_X1 port map( A1 => a(9), A2 => n6, B1 => c(9), B2 => n7, ZN => n2
                           );
   U8 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => y(8));
   U9 : AOI22_X1 port map( A1 => d(8), A2 => n1, B1 => b(8), B2 => n5, ZN => n9
                           );
   U10 : AOI22_X1 port map( A1 => a(8), A2 => n6, B1 => c(8), B2 => n7, ZN => 
                           n8);
   U11 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => y(7));
   U12 : AOI22_X1 port map( A1 => d(7), A2 => n1, B1 => b(7), B2 => n5, ZN => 
                           n11);
   U13 : AOI22_X1 port map( A1 => a(7), A2 => n6, B1 => c(7), B2 => n7, ZN => 
                           n10);
   U14 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => y(6));
   U15 : AOI22_X1 port map( A1 => d(6), A2 => n1, B1 => b(6), B2 => n5, ZN => 
                           n13);
   U16 : AOI22_X1 port map( A1 => a(6), A2 => n6, B1 => c(6), B2 => n7, ZN => 
                           n12);
   U17 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => y(5));
   U18 : AOI22_X1 port map( A1 => d(5), A2 => n1, B1 => b(5), B2 => n5, ZN => 
                           n15);
   U19 : AOI22_X1 port map( A1 => a(5), A2 => n6, B1 => c(5), B2 => n7, ZN => 
                           n14);
   U20 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => y(4));
   U21 : AOI22_X1 port map( A1 => d(4), A2 => n1, B1 => b(4), B2 => n5, ZN => 
                           n17);
   U22 : AOI22_X1 port map( A1 => a(4), A2 => n6, B1 => c(4), B2 => n7, ZN => 
                           n16);
   U23 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => y(3));
   U24 : AOI22_X1 port map( A1 => d(3), A2 => n1, B1 => b(3), B2 => n5, ZN => 
                           n19);
   U25 : AOI22_X1 port map( A1 => a(3), A2 => n6, B1 => c(3), B2 => n7, ZN => 
                           n18);
   U26 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => y(39));
   U27 : AOI22_X1 port map( A1 => d(39), A2 => n1, B1 => b(39), B2 => n5, ZN =>
                           n21);
   U28 : AOI22_X1 port map( A1 => a(39), A2 => n6, B1 => c(39), B2 => n7, ZN =>
                           n20);
   U29 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => y(38));
   U30 : AOI22_X1 port map( A1 => d(38), A2 => n1, B1 => b(38), B2 => n5, ZN =>
                           n23);
   U31 : AOI22_X1 port map( A1 => a(38), A2 => n6, B1 => c(38), B2 => n7, ZN =>
                           n22);
   U32 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => y(37));
   U33 : AOI22_X1 port map( A1 => d(37), A2 => n1, B1 => b(37), B2 => n5, ZN =>
                           n25);
   U34 : AOI22_X1 port map( A1 => a(37), A2 => n6, B1 => c(37), B2 => n7, ZN =>
                           n24);
   U35 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => y(36));
   U36 : AOI22_X1 port map( A1 => d(36), A2 => n1, B1 => b(36), B2 => n5, ZN =>
                           n27);
   U37 : AOI22_X1 port map( A1 => a(36), A2 => n6, B1 => c(36), B2 => n7, ZN =>
                           n26);
   U38 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => y(35));
   U39 : AOI22_X1 port map( A1 => d(35), A2 => n1, B1 => b(35), B2 => n5, ZN =>
                           n29);
   U40 : AOI22_X1 port map( A1 => a(35), A2 => n6, B1 => c(35), B2 => n7, ZN =>
                           n28);
   U41 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => y(34));
   U42 : AOI22_X1 port map( A1 => d(34), A2 => n1, B1 => b(34), B2 => n5, ZN =>
                           n31);
   U43 : AOI22_X1 port map( A1 => a(34), A2 => n6, B1 => c(34), B2 => n7, ZN =>
                           n30);
   U44 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => y(33));
   U45 : AOI22_X1 port map( A1 => d(33), A2 => n1, B1 => b(33), B2 => n5, ZN =>
                           n33);
   U46 : AOI22_X1 port map( A1 => a(33), A2 => n6, B1 => c(33), B2 => n7, ZN =>
                           n32);
   U47 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => y(32));
   U48 : AOI22_X1 port map( A1 => d(32), A2 => n1, B1 => b(32), B2 => n5, ZN =>
                           n35);
   U49 : AOI22_X1 port map( A1 => a(32), A2 => n6, B1 => c(32), B2 => n7, ZN =>
                           n34);
   U50 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => y(31));
   U51 : AOI22_X1 port map( A1 => d(31), A2 => n1, B1 => b(31), B2 => n5, ZN =>
                           n37);
   U52 : AOI22_X1 port map( A1 => a(31), A2 => n6, B1 => c(31), B2 => n7, ZN =>
                           n36);
   U53 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => y(30));
   U54 : AOI22_X1 port map( A1 => d(30), A2 => n1, B1 => b(30), B2 => n5, ZN =>
                           n39);
   U55 : AOI22_X1 port map( A1 => a(30), A2 => n6, B1 => c(30), B2 => n7, ZN =>
                           n38);
   U56 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => y(2));
   U57 : AOI22_X1 port map( A1 => d(2), A2 => n1, B1 => b(2), B2 => n5, ZN => 
                           n41);
   U58 : AOI22_X1 port map( A1 => a(2), A2 => n6, B1 => c(2), B2 => n7, ZN => 
                           n40);
   U59 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => y(29));
   U60 : AOI22_X1 port map( A1 => d(29), A2 => n1, B1 => b(29), B2 => n5, ZN =>
                           n43);
   U61 : AOI22_X1 port map( A1 => a(29), A2 => n6, B1 => c(29), B2 => n7, ZN =>
                           n42);
   U62 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => y(28));
   U63 : AOI22_X1 port map( A1 => d(28), A2 => n1, B1 => b(28), B2 => n5, ZN =>
                           n45);
   U64 : AOI22_X1 port map( A1 => a(28), A2 => n6, B1 => c(28), B2 => n7, ZN =>
                           n44);
   U65 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => y(27));
   U66 : AOI22_X1 port map( A1 => d(27), A2 => n1, B1 => b(27), B2 => n5, ZN =>
                           n47);
   U67 : AOI22_X1 port map( A1 => a(27), A2 => n6, B1 => c(27), B2 => n7, ZN =>
                           n46);
   U68 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => y(26));
   U69 : AOI22_X1 port map( A1 => d(26), A2 => n1, B1 => b(26), B2 => n5, ZN =>
                           n49);
   U70 : AOI22_X1 port map( A1 => a(26), A2 => n6, B1 => c(26), B2 => n7, ZN =>
                           n48);
   U71 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => y(25));
   U72 : AOI22_X1 port map( A1 => d(25), A2 => n1, B1 => b(25), B2 => n5, ZN =>
                           n51);
   U73 : AOI22_X1 port map( A1 => a(25), A2 => n6, B1 => c(25), B2 => n7, ZN =>
                           n50);
   U74 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => y(24));
   U75 : AOI22_X1 port map( A1 => d(24), A2 => n1, B1 => b(24), B2 => n5, ZN =>
                           n53);
   U76 : AOI22_X1 port map( A1 => a(24), A2 => n6, B1 => c(24), B2 => n7, ZN =>
                           n52);
   U77 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => y(23));
   U78 : AOI22_X1 port map( A1 => d(23), A2 => n1, B1 => b(23), B2 => n5, ZN =>
                           n55);
   U79 : AOI22_X1 port map( A1 => a(23), A2 => n6, B1 => c(23), B2 => n7, ZN =>
                           n54);
   U80 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => y(22));
   U81 : AOI22_X1 port map( A1 => d(22), A2 => n1, B1 => b(22), B2 => n5, ZN =>
                           n57);
   U82 : AOI22_X1 port map( A1 => a(22), A2 => n6, B1 => c(22), B2 => n7, ZN =>
                           n56);
   U83 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => y(21));
   U84 : AOI22_X1 port map( A1 => d(21), A2 => n1, B1 => b(21), B2 => n5, ZN =>
                           n59);
   U85 : AOI22_X1 port map( A1 => a(21), A2 => n6, B1 => c(21), B2 => n7, ZN =>
                           n58);
   U86 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => y(20));
   U87 : AOI22_X1 port map( A1 => d(20), A2 => n1, B1 => b(20), B2 => n5, ZN =>
                           n61);
   U88 : AOI22_X1 port map( A1 => a(20), A2 => n6, B1 => c(20), B2 => n7, ZN =>
                           n60);
   U89 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => y(1));
   U90 : AOI22_X1 port map( A1 => d(1), A2 => n1, B1 => b(1), B2 => n5, ZN => 
                           n63);
   U91 : AOI22_X1 port map( A1 => a(1), A2 => n6, B1 => c(1), B2 => n7, ZN => 
                           n62);
   U92 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => y(19));
   U93 : AOI22_X1 port map( A1 => d(19), A2 => n1, B1 => b(19), B2 => n5, ZN =>
                           n65);
   U94 : AOI22_X1 port map( A1 => a(19), A2 => n6, B1 => c(19), B2 => n7, ZN =>
                           n64);
   U95 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => y(18));
   U96 : AOI22_X1 port map( A1 => d(18), A2 => n1, B1 => b(18), B2 => n5, ZN =>
                           n67);
   U97 : AOI22_X1 port map( A1 => a(18), A2 => n6, B1 => c(18), B2 => n7, ZN =>
                           n66);
   U98 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => y(17));
   U99 : AOI22_X1 port map( A1 => d(17), A2 => n1, B1 => b(17), B2 => n5, ZN =>
                           n69);
   U100 : AOI22_X1 port map( A1 => a(17), A2 => n6, B1 => c(17), B2 => n7, ZN 
                           => n68);
   U101 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => y(16));
   U102 : AOI22_X1 port map( A1 => d(16), A2 => n1, B1 => b(16), B2 => n5, ZN 
                           => n71);
   U103 : AOI22_X1 port map( A1 => a(16), A2 => n6, B1 => c(16), B2 => n7, ZN 
                           => n70);
   U104 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => y(15));
   U105 : AOI22_X1 port map( A1 => d(15), A2 => n1, B1 => b(15), B2 => n5, ZN 
                           => n73);
   U106 : AOI22_X1 port map( A1 => a(15), A2 => n6, B1 => c(15), B2 => n7, ZN 
                           => n72);
   U107 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => y(14));
   U108 : AOI22_X1 port map( A1 => d(14), A2 => n1, B1 => b(14), B2 => n5, ZN 
                           => n75);
   U109 : AOI22_X1 port map( A1 => a(14), A2 => n6, B1 => c(14), B2 => n7, ZN 
                           => n74);
   U110 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => y(13));
   U111 : AOI22_X1 port map( A1 => d(13), A2 => n1, B1 => b(13), B2 => n5, ZN 
                           => n77);
   U112 : AOI22_X1 port map( A1 => a(13), A2 => n6, B1 => c(13), B2 => n7, ZN 
                           => n76);
   U113 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => y(12));
   U114 : AOI22_X1 port map( A1 => d(12), A2 => n1, B1 => b(12), B2 => n5, ZN 
                           => n79);
   U115 : AOI22_X1 port map( A1 => a(12), A2 => n6, B1 => c(12), B2 => n7, ZN 
                           => n78);
   U116 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => y(11));
   U117 : AOI22_X1 port map( A1 => d(11), A2 => n1, B1 => b(11), B2 => n5, ZN 
                           => n81);
   U118 : AOI22_X1 port map( A1 => a(11), A2 => n6, B1 => c(11), B2 => n7, ZN 
                           => n80);
   U119 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => y(10));
   U120 : AOI22_X1 port map( A1 => d(10), A2 => n1, B1 => b(10), B2 => n5, ZN 
                           => n83);
   U121 : AOI22_X1 port map( A1 => a(10), A2 => n6, B1 => c(10), B2 => n7, ZN 
                           => n82);
   U122 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => y(0));
   U123 : AOI22_X1 port map( A1 => d(0), A2 => n1, B1 => b(0), B2 => n5, ZN => 
                           n85);
   U124 : NOR3_X1 port map( A1 => n6, A2 => n7, A3 => n5, ZN => n4);
   U125 : AOI22_X1 port map( A1 => a(0), A2 => n6, B1 => c(0), B2 => n7, ZN => 
                           n84);
   U126 : INV_X1 port map( A => sel(1), ZN => n86);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N40_0 is

   port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (39 downto 0));

end MUX21_N40_0;

architecture SYN_beh of MUX21_N40_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));
   U2 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U3 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U4 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U5 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U6 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U7 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U8 : MUX2_X1 port map( A => a(39), B => b(39), S => sel, Z => y(39));
   U9 : MUX2_X1 port map( A => a(38), B => b(38), S => sel, Z => y(38));
   U10 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U11 : MUX2_X1 port map( A => a(32), B => b(32), S => sel, Z => y(32));
   U12 : MUX2_X1 port map( A => a(33), B => b(33), S => sel, Z => y(33));
   U13 : MUX2_X1 port map( A => a(34), B => b(34), S => sel, Z => y(34));
   U14 : MUX2_X1 port map( A => a(35), B => b(35), S => sel, Z => y(35));
   U15 : MUX2_X1 port map( A => a(36), B => b(36), S => sel, Z => y(36));
   U16 : MUX2_X1 port map( A => a(37), B => b(37), S => sel, Z => y(37));
   U17 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U18 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U19 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U20 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U21 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U22 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U23 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U24 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U25 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U26 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U27 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U28 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U29 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U30 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U31 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U32 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U33 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U34 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U35 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U36 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U37 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U38 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U39 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U40 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT7 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT7;

architecture SYN_behavioral of shift_NBIT32_SHIFT7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_2a_31_port, neg_2a_30_port, n3, n4, n5, n6, n7, n8
      , n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_16_port, neg_2a_20_port, 
      neg_2a_24_port, neg_2a_27_port, neg_2a_17_port, neg_2a_19_port, 
      neg_2a_23_port, neg_2a_26_port, neg_2a_18_port, neg_2a_22_port, 
      neg_2a_25_port, neg_2a_29_port, neg_2a_21_port, neg_2a_28_port, n31, n32,
      n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47
      : std_logic;

begin
   pos_a <= ( a(15), a(15), a(15), a(14), a(13), a(12), a(11), a(10), a(9), 
      a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   neg_a <= ( neg_2a_31_port, neg_2a_31_port, neg_2a_30_port, neg_2a_29_port, 
      neg_2a_28_port, neg_2a_27_port, neg_2a_26_port, neg_2a_25_port, 
      neg_2a_24_port, neg_2a_23_port, neg_2a_22_port, neg_2a_21_port, 
      neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, 
      neg_2a_16_port, a(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   pos_2a <= ( a(15), a(15), a(14), a(13), a(12), a(11), a(10), a(9), a(8), 
      a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   neg_2a <= ( neg_2a_31_port, neg_2a_30_port, neg_2a_29_port, neg_2a_28_port, 
      neg_2a_27_port, neg_2a_26_port, neg_2a_25_port, neg_2a_24_port, 
      neg_2a_23_port, neg_2a_22_port, neg_2a_21_port, neg_2a_20_port, 
      neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, neg_2a_16_port, a(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : XNOR2_X1 port map( A => n31, B => n32, ZN => neg_2a_31_port);
   U3 : NAND2_X1 port map( A1 => n31, A2 => n16, ZN => n32);
   U4 : XOR2_X1 port map( A => n31, B => n16, Z => neg_2a_30_port);
   U5 : AND2_X1 port map( A1 => n34, A2 => n33, ZN => n3);
   U6 : AND2_X1 port map( A1 => n41, A2 => n11, ZN => n4);
   U7 : AND2_X1 port map( A1 => n42, A2 => n4, ZN => n5);
   U8 : AND2_X1 port map( A1 => n35, A2 => n3, ZN => n6);
   U9 : AND2_X1 port map( A1 => n36, A2 => n6, ZN => n7);
   U10 : AND2_X1 port map( A1 => n37, A2 => n7, ZN => n8);
   U11 : AND2_X1 port map( A1 => n38, A2 => n8, ZN => n9);
   U12 : AND2_X1 port map( A1 => n39, A2 => n9, ZN => n10);
   U13 : AND2_X1 port map( A1 => n40, A2 => n10, ZN => n11);
   U14 : AND2_X1 port map( A1 => n43, A2 => n5, ZN => n12);
   U15 : AND2_X1 port map( A1 => n44, A2 => n12, ZN => n13);
   U16 : AND2_X1 port map( A1 => n45, A2 => n13, ZN => n14);
   U17 : AND2_X1 port map( A1 => n46, A2 => n14, ZN => n15);
   U18 : AND2_X1 port map( A1 => n47, A2 => n15, ZN => n16);
   U19 : XOR2_X1 port map( A => n34, B => n33, Z => neg_2a_16_port);
   U20 : XOR2_X1 port map( A => n38, B => n8, Z => neg_2a_20_port);
   U21 : XOR2_X1 port map( A => n42, B => n4, Z => neg_2a_24_port);
   U22 : XOR2_X1 port map( A => n45, B => n13, Z => neg_2a_27_port);
   U23 : XOR2_X1 port map( A => n35, B => n3, Z => neg_2a_17_port);
   U24 : XOR2_X1 port map( A => n37, B => n7, Z => neg_2a_19_port);
   U25 : XOR2_X1 port map( A => n41, B => n11, Z => neg_2a_23_port);
   U26 : XOR2_X1 port map( A => n44, B => n12, Z => neg_2a_26_port);
   U27 : XOR2_X1 port map( A => n36, B => n6, Z => neg_2a_18_port);
   U28 : XOR2_X1 port map( A => n40, B => n10, Z => neg_2a_22_port);
   U29 : XOR2_X1 port map( A => n43, B => n5, Z => neg_2a_25_port);
   U30 : XOR2_X1 port map( A => n47, B => n15, Z => neg_2a_29_port);
   U31 : XOR2_X1 port map( A => n39, B => n9, Z => neg_2a_21_port);
   U32 : XOR2_X1 port map( A => n46, B => n14, Z => neg_2a_28_port);
   U33 : INV_X1 port map( A => a(15), ZN => n31);
   U34 : INV_X1 port map( A => a(14), ZN => n47);
   U35 : INV_X1 port map( A => a(13), ZN => n46);
   U36 : INV_X1 port map( A => a(12), ZN => n45);
   U37 : INV_X1 port map( A => a(11), ZN => n44);
   U38 : INV_X1 port map( A => a(10), ZN => n43);
   U39 : INV_X1 port map( A => a(9), ZN => n42);
   U40 : INV_X1 port map( A => a(8), ZN => n41);
   U41 : INV_X1 port map( A => a(7), ZN => n40);
   U42 : INV_X1 port map( A => a(6), ZN => n39);
   U43 : INV_X1 port map( A => a(5), ZN => n38);
   U44 : INV_X1 port map( A => a(4), ZN => n37);
   U45 : INV_X1 port map( A => a(3), ZN => n36);
   U46 : INV_X1 port map( A => a(2), ZN => n35);
   U47 : INV_X1 port map( A => a(1), ZN => n34);
   U48 : INV_X1 port map( A => a(0), ZN => n33);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT6 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT6;

architecture SYN_behavioral of shift_NBIT32_SHIFT6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_2a_29_port, neg_2a_28_port, n3, n4, n5, n6, n7, n8
      , n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_14_port, neg_2a_18_port, 
      neg_2a_22_port, neg_2a_25_port, neg_2a_15_port, neg_2a_17_port, 
      neg_2a_21_port, neg_2a_24_port, neg_2a_16_port, neg_2a_20_port, 
      neg_2a_23_port, neg_2a_27_port, neg_2a_19_port, neg_2a_26_port, n31, n32,
      n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47
      : std_logic;

begin
   pos_a <= ( a(15), a(15), a(15), a(15), a(15), a(14), a(13), a(12), a(11), 
      a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   neg_a <= ( neg_2a_29_port, neg_2a_29_port, neg_2a_29_port, neg_2a_29_port, 
      neg_2a_28_port, neg_2a_27_port, neg_2a_26_port, neg_2a_25_port, 
      neg_2a_24_port, neg_2a_23_port, neg_2a_22_port, neg_2a_21_port, 
      neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, 
      neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   pos_2a <= ( a(15), a(15), a(15), a(15), a(14), a(13), a(12), a(11), a(10), 
      a(9), a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   neg_2a <= ( neg_2a_29_port, neg_2a_29_port, neg_2a_29_port, neg_2a_28_port, 
      neg_2a_27_port, neg_2a_26_port, neg_2a_25_port, neg_2a_24_port, 
      neg_2a_23_port, neg_2a_22_port, neg_2a_21_port, neg_2a_20_port, 
      neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, neg_2a_16_port, 
      neg_2a_15_port, neg_2a_14_port, a(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : XNOR2_X1 port map( A => n31, B => n32, ZN => neg_2a_29_port);
   U3 : NAND2_X1 port map( A1 => n31, A2 => n16, ZN => n32);
   U4 : XOR2_X1 port map( A => n31, B => n16, Z => neg_2a_28_port);
   U5 : AND2_X1 port map( A1 => n34, A2 => n33, ZN => n3);
   U6 : AND2_X1 port map( A1 => n38, A2 => n8, ZN => n4);
   U7 : AND2_X1 port map( A1 => n45, A2 => n14, ZN => n5);
   U8 : AND2_X1 port map( A1 => n35, A2 => n3, ZN => n6);
   U9 : AND2_X1 port map( A1 => n36, A2 => n6, ZN => n7);
   U10 : AND2_X1 port map( A1 => n37, A2 => n7, ZN => n8);
   U11 : AND2_X1 port map( A1 => n39, A2 => n4, ZN => n9);
   U12 : AND2_X1 port map( A1 => n40, A2 => n9, ZN => n10);
   U13 : AND2_X1 port map( A1 => n41, A2 => n10, ZN => n11);
   U14 : AND2_X1 port map( A1 => n42, A2 => n11, ZN => n12);
   U15 : AND2_X1 port map( A1 => n43, A2 => n12, ZN => n13);
   U16 : AND2_X1 port map( A1 => n44, A2 => n13, ZN => n14);
   U17 : AND2_X1 port map( A1 => n46, A2 => n5, ZN => n15);
   U18 : AND2_X1 port map( A1 => n47, A2 => n15, ZN => n16);
   U19 : XOR2_X1 port map( A => n34, B => n33, Z => neg_2a_14_port);
   U20 : XOR2_X1 port map( A => n38, B => n8, Z => neg_2a_18_port);
   U21 : XOR2_X1 port map( A => n42, B => n11, Z => neg_2a_22_port);
   U22 : XOR2_X1 port map( A => n45, B => n14, Z => neg_2a_25_port);
   U23 : XOR2_X1 port map( A => n35, B => n3, Z => neg_2a_15_port);
   U24 : XOR2_X1 port map( A => n37, B => n7, Z => neg_2a_17_port);
   U25 : XOR2_X1 port map( A => n41, B => n10, Z => neg_2a_21_port);
   U26 : XOR2_X1 port map( A => n44, B => n13, Z => neg_2a_24_port);
   U27 : XOR2_X1 port map( A => n36, B => n6, Z => neg_2a_16_port);
   U28 : XOR2_X1 port map( A => n40, B => n9, Z => neg_2a_20_port);
   U29 : XOR2_X1 port map( A => n43, B => n12, Z => neg_2a_23_port);
   U30 : XOR2_X1 port map( A => n47, B => n15, Z => neg_2a_27_port);
   U31 : XOR2_X1 port map( A => n39, B => n4, Z => neg_2a_19_port);
   U32 : XOR2_X1 port map( A => n46, B => n5, Z => neg_2a_26_port);
   U33 : INV_X1 port map( A => a(15), ZN => n31);
   U34 : INV_X1 port map( A => a(14), ZN => n47);
   U35 : INV_X1 port map( A => a(13), ZN => n46);
   U36 : INV_X1 port map( A => a(12), ZN => n45);
   U37 : INV_X1 port map( A => a(11), ZN => n44);
   U38 : INV_X1 port map( A => a(10), ZN => n43);
   U39 : INV_X1 port map( A => a(9), ZN => n42);
   U40 : INV_X1 port map( A => a(8), ZN => n41);
   U41 : INV_X1 port map( A => a(7), ZN => n40);
   U42 : INV_X1 port map( A => a(6), ZN => n39);
   U43 : INV_X1 port map( A => a(5), ZN => n38);
   U44 : INV_X1 port map( A => a(4), ZN => n37);
   U45 : INV_X1 port map( A => a(3), ZN => n36);
   U46 : INV_X1 port map( A => a(2), ZN => n35);
   U47 : INV_X1 port map( A => a(1), ZN => n34);
   U48 : INV_X1 port map( A => a(0), ZN => n33);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT5 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT5;

architecture SYN_behavioral of shift_NBIT32_SHIFT5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_2a_27_port, neg_2a_26_port, n3, n4, n5, n6, n7, n8
      , n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_12_port, neg_2a_16_port, 
      neg_2a_20_port, neg_2a_23_port, neg_2a_13_port, neg_2a_15_port, 
      neg_2a_19_port, neg_2a_22_port, neg_2a_14_port, neg_2a_18_port, 
      neg_2a_21_port, neg_2a_25_port, neg_2a_17_port, neg_2a_24_port, 
      pos_2a_26_port, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48 : std_logic;

begin
   pos_a <= ( pos_2a_26_port, pos_2a_26_port, pos_2a_26_port, pos_2a_26_port, 
      pos_2a_26_port, pos_2a_26_port, pos_2a_26_port, a(14), a(13), a(12), 
      a(11), a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0),
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port );
   neg_a <= ( neg_2a_27_port, neg_2a_27_port, neg_2a_27_port, neg_2a_27_port, 
      neg_2a_27_port, neg_2a_27_port, neg_2a_26_port, neg_2a_25_port, 
      neg_2a_24_port, neg_2a_23_port, neg_2a_22_port, neg_2a_21_port, 
      neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, 
      neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, neg_2a_13_port, 
      neg_2a_12_port, a(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port );
   pos_2a <= ( pos_2a_26_port, pos_2a_26_port, pos_2a_26_port, pos_2a_26_port, 
      pos_2a_26_port, pos_2a_26_port, a(14), a(13), a(12), a(11), a(10), a(9), 
      a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port );
   neg_2a <= ( neg_2a_27_port, neg_2a_27_port, neg_2a_27_port, neg_2a_27_port, 
      neg_2a_27_port, neg_2a_26_port, neg_2a_25_port, neg_2a_24_port, 
      neg_2a_23_port, neg_2a_22_port, neg_2a_21_port, neg_2a_20_port, 
      neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, neg_2a_16_port, 
      neg_2a_15_port, neg_2a_14_port, neg_2a_13_port, neg_2a_12_port, a(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : XNOR2_X1 port map( A => n32, B => n33, ZN => neg_2a_27_port);
   U3 : NAND2_X1 port map( A1 => n32, A2 => n16, ZN => n33);
   U4 : XOR2_X1 port map( A => n32, B => n16, Z => neg_2a_26_port);
   U5 : INV_X1 port map( A => a(15), ZN => n32);
   U6 : AND2_X1 port map( A1 => n35, A2 => n34, ZN => n3);
   U7 : AND2_X1 port map( A1 => n39, A2 => n8, ZN => n4);
   U8 : AND2_X1 port map( A1 => n36, A2 => n3, ZN => n5);
   U9 : AND2_X1 port map( A1 => n43, A2 => n11, ZN => n6);
   U10 : AND2_X1 port map( A1 => n37, A2 => n5, ZN => n7);
   U11 : AND2_X1 port map( A1 => n38, A2 => n7, ZN => n8);
   U12 : AND2_X1 port map( A1 => n40, A2 => n4, ZN => n9);
   U13 : AND2_X1 port map( A1 => n41, A2 => n9, ZN => n10);
   U14 : AND2_X1 port map( A1 => n42, A2 => n10, ZN => n11);
   U15 : AND2_X1 port map( A1 => n44, A2 => n6, ZN => n12);
   U16 : AND2_X1 port map( A1 => n45, A2 => n12, ZN => n13);
   U17 : AND2_X1 port map( A1 => n46, A2 => n13, ZN => n14);
   U18 : AND2_X1 port map( A1 => n47, A2 => n14, ZN => n15);
   U19 : AND2_X1 port map( A1 => n48, A2 => n15, ZN => n16);
   U20 : XOR2_X1 port map( A => n35, B => n34, Z => neg_2a_12_port);
   U21 : XOR2_X1 port map( A => n39, B => n8, Z => neg_2a_16_port);
   U22 : XOR2_X1 port map( A => n43, B => n11, Z => neg_2a_20_port);
   U23 : XOR2_X1 port map( A => n46, B => n13, Z => neg_2a_23_port);
   U24 : XOR2_X1 port map( A => n36, B => n3, Z => neg_2a_13_port);
   U25 : XOR2_X1 port map( A => n38, B => n7, Z => neg_2a_15_port);
   U26 : XOR2_X1 port map( A => n42, B => n10, Z => neg_2a_19_port);
   U27 : XOR2_X1 port map( A => n45, B => n12, Z => neg_2a_22_port);
   U28 : XOR2_X1 port map( A => n37, B => n5, Z => neg_2a_14_port);
   U29 : XOR2_X1 port map( A => n41, B => n9, Z => neg_2a_18_port);
   U30 : XOR2_X1 port map( A => n44, B => n6, Z => neg_2a_21_port);
   U31 : XOR2_X1 port map( A => n48, B => n15, Z => neg_2a_25_port);
   U32 : XOR2_X1 port map( A => n40, B => n4, Z => neg_2a_17_port);
   U33 : XOR2_X1 port map( A => n47, B => n14, Z => neg_2a_24_port);
   U34 : INV_X1 port map( A => n32, ZN => pos_2a_26_port);
   U35 : INV_X1 port map( A => a(14), ZN => n48);
   U36 : INV_X1 port map( A => a(13), ZN => n47);
   U37 : INV_X1 port map( A => a(12), ZN => n46);
   U38 : INV_X1 port map( A => a(11), ZN => n45);
   U39 : INV_X1 port map( A => a(10), ZN => n44);
   U40 : INV_X1 port map( A => a(9), ZN => n43);
   U41 : INV_X1 port map( A => a(8), ZN => n42);
   U42 : INV_X1 port map( A => a(7), ZN => n41);
   U43 : INV_X1 port map( A => a(6), ZN => n40);
   U44 : INV_X1 port map( A => a(5), ZN => n39);
   U45 : INV_X1 port map( A => a(4), ZN => n38);
   U46 : INV_X1 port map( A => a(3), ZN => n37);
   U47 : INV_X1 port map( A => a(2), ZN => n36);
   U48 : INV_X1 port map( A => a(1), ZN => n35);
   U49 : INV_X1 port map( A => a(0), ZN => n34);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT4 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT4;

architecture SYN_behavioral of shift_NBIT32_SHIFT4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_a_31, n1, neg_2a_24_port, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_10_port, neg_2a_14_port, 
      neg_2a_18_port, neg_2a_21_port, neg_2a_11_port, neg_2a_13_port, 
      neg_2a_17_port, neg_2a_20_port, neg_2a_12_port, neg_2a_16_port, 
      neg_2a_19_port, neg_2a_23_port, neg_2a_15_port, neg_2a_22_port, 
      pos_2a_24_port, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48 : std_logic;

begin
   pos_a <= ( pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, 
      pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, 
      pos_2a_24_port, a(14), a(13), a(12), a(11), a(10), a(9), a(8), a(7), a(6)
      , a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port );
   neg_a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_2a_24_port, neg_2a_23_port, neg_2a_22_port, 
      neg_2a_21_port, neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, 
      neg_2a_17_port, neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, 
      neg_2a_13_port, neg_2a_12_port, neg_2a_11_port, neg_2a_10_port, a(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   pos_2a <= ( pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, 
      pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, pos_2a_24_port, a(14), 
      a(13), a(12), a(11), a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), 
      a(2), a(1), a(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port );
   neg_2a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_2a_24_port, neg_2a_23_port, neg_2a_22_port, neg_2a_21_port,
      neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, 
      neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, neg_2a_13_port, 
      neg_2a_12_port, neg_2a_11_port, neg_2a_10_port, a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND2_X1 port map( A1 => n32, A2 => n16, ZN => n1);
   U3 : INV_X1 port map( A => n33, ZN => neg_a_31);
   U4 : XNOR2_X1 port map( A => n32, B => n1, ZN => n33);
   U5 : XOR2_X1 port map( A => n32, B => n16, Z => neg_2a_24_port);
   U6 : INV_X1 port map( A => a(15), ZN => n32);
   U7 : AND2_X1 port map( A1 => n35, A2 => n34, ZN => n3);
   U8 : AND2_X1 port map( A1 => n39, A2 => n7, ZN => n4);
   U9 : AND2_X1 port map( A1 => n36, A2 => n3, ZN => n5);
   U10 : AND2_X1 port map( A1 => n37, A2 => n5, ZN => n6);
   U11 : AND2_X1 port map( A1 => n38, A2 => n6, ZN => n7);
   U12 : AND2_X1 port map( A1 => n41, A2 => n10, ZN => n8);
   U13 : AND2_X1 port map( A1 => n46, A2 => n14, ZN => n9);
   U14 : AND2_X1 port map( A1 => n40, A2 => n4, ZN => n10);
   U15 : AND2_X1 port map( A1 => n42, A2 => n8, ZN => n11);
   U16 : AND2_X1 port map( A1 => n43, A2 => n11, ZN => n12);
   U17 : AND2_X1 port map( A1 => n44, A2 => n12, ZN => n13);
   U18 : AND2_X1 port map( A1 => n45, A2 => n13, ZN => n14);
   U19 : AND2_X1 port map( A1 => n47, A2 => n9, ZN => n15);
   U20 : AND2_X1 port map( A1 => n48, A2 => n15, ZN => n16);
   U21 : XOR2_X1 port map( A => n35, B => n34, Z => neg_2a_10_port);
   U22 : XOR2_X1 port map( A => n39, B => n7, Z => neg_2a_14_port);
   U23 : XOR2_X1 port map( A => n43, B => n11, Z => neg_2a_18_port);
   U24 : XOR2_X1 port map( A => n46, B => n14, Z => neg_2a_21_port);
   U25 : XOR2_X1 port map( A => n36, B => n3, Z => neg_2a_11_port);
   U26 : XOR2_X1 port map( A => n38, B => n6, Z => neg_2a_13_port);
   U27 : XOR2_X1 port map( A => n42, B => n8, Z => neg_2a_17_port);
   U28 : XOR2_X1 port map( A => n45, B => n13, Z => neg_2a_20_port);
   U29 : XOR2_X1 port map( A => n37, B => n5, Z => neg_2a_12_port);
   U30 : XOR2_X1 port map( A => n41, B => n10, Z => neg_2a_16_port);
   U31 : XOR2_X1 port map( A => n44, B => n12, Z => neg_2a_19_port);
   U32 : XOR2_X1 port map( A => n48, B => n15, Z => neg_2a_23_port);
   U33 : XOR2_X1 port map( A => n40, B => n4, Z => neg_2a_15_port);
   U34 : XOR2_X1 port map( A => n47, B => n9, Z => neg_2a_22_port);
   U35 : INV_X1 port map( A => n32, ZN => pos_2a_24_port);
   U36 : INV_X1 port map( A => a(14), ZN => n48);
   U37 : INV_X1 port map( A => a(13), ZN => n47);
   U38 : INV_X1 port map( A => a(12), ZN => n46);
   U39 : INV_X1 port map( A => a(11), ZN => n45);
   U40 : INV_X1 port map( A => a(10), ZN => n44);
   U41 : INV_X1 port map( A => a(9), ZN => n43);
   U42 : INV_X1 port map( A => a(8), ZN => n42);
   U43 : INV_X1 port map( A => a(7), ZN => n41);
   U44 : INV_X1 port map( A => a(6), ZN => n40);
   U45 : INV_X1 port map( A => a(5), ZN => n39);
   U46 : INV_X1 port map( A => a(4), ZN => n38);
   U47 : INV_X1 port map( A => a(3), ZN => n37);
   U48 : INV_X1 port map( A => a(2), ZN => n36);
   U49 : INV_X1 port map( A => a(1), ZN => n35);
   U50 : INV_X1 port map( A => a(0), ZN => n34);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT3 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT3;

architecture SYN_behavioral of shift_NBIT32_SHIFT3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_a_31, n1, neg_2a_22_port, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_8_port, neg_2a_12_port, 
      neg_2a_16_port, neg_2a_19_port, neg_2a_9_port, neg_2a_11_port, 
      neg_2a_15_port, neg_2a_18_port, neg_2a_10_port, neg_2a_14_port, 
      neg_2a_17_port, neg_2a_21_port, neg_2a_13_port, neg_2a_20_port, 
      pos_2a_22_port, pos_a_23_port, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49 : std_logic;

begin
   pos_a <= ( pos_a_23_port, pos_a_23_port, pos_a_23_port, pos_a_23_port, 
      pos_a_23_port, pos_a_23_port, pos_a_23_port, pos_a_23_port, pos_a_23_port
      , pos_2a_22_port, pos_2a_22_port, a(14), a(13), a(12), a(11), a(10), a(9)
      , a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   neg_a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_2a_22_port, neg_2a_21_port, 
      neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, 
      neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, neg_2a_13_port, 
      neg_2a_12_port, neg_2a_11_port, neg_2a_10_port, neg_2a_9_port, 
      neg_2a_8_port, a(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   pos_2a <= ( pos_2a_22_port, pos_2a_22_port, pos_2a_22_port, pos_2a_22_port, 
      pos_2a_22_port, pos_2a_22_port, pos_2a_22_port, pos_2a_22_port, 
      pos_2a_22_port, pos_2a_22_port, a(14), a(13), a(12), a(11), a(10), a(9), 
      a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port );
   neg_2a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_2a_22_port, neg_2a_21_port, 
      neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, 
      neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, neg_2a_13_port, 
      neg_2a_12_port, neg_2a_11_port, neg_2a_10_port, neg_2a_9_port, 
      neg_2a_8_port, a(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND2_X1 port map( A1 => n33, A2 => n16, ZN => n1);
   U3 : INV_X1 port map( A => n34, ZN => neg_a_31);
   U4 : XNOR2_X1 port map( A => n33, B => n1, ZN => n34);
   U5 : XOR2_X1 port map( A => n33, B => n16, Z => neg_2a_22_port);
   U6 : INV_X1 port map( A => a(15), ZN => n33);
   U7 : AND2_X1 port map( A1 => n36, A2 => n35, ZN => n3);
   U8 : AND2_X1 port map( A1 => n40, A2 => n6, ZN => n4);
   U9 : AND2_X1 port map( A1 => n37, A2 => n3, ZN => n5);
   U10 : AND2_X1 port map( A1 => n39, A2 => n7, ZN => n6);
   U11 : AND2_X1 port map( A1 => n38, A2 => n5, ZN => n7);
   U12 : AND2_X1 port map( A1 => n41, A2 => n4, ZN => n8);
   U13 : AND2_X1 port map( A1 => n42, A2 => n8, ZN => n9);
   U14 : AND2_X1 port map( A1 => n43, A2 => n9, ZN => n10);
   U15 : AND2_X1 port map( A1 => n44, A2 => n10, ZN => n11);
   U16 : AND2_X1 port map( A1 => n46, A2 => n13, ZN => n12);
   U17 : AND2_X1 port map( A1 => n45, A2 => n11, ZN => n13);
   U18 : AND2_X1 port map( A1 => n47, A2 => n12, ZN => n14);
   U19 : AND2_X1 port map( A1 => n48, A2 => n14, ZN => n15);
   U20 : AND2_X1 port map( A1 => n49, A2 => n15, ZN => n16);
   U21 : XOR2_X1 port map( A => n36, B => n35, Z => neg_2a_8_port);
   U22 : XOR2_X1 port map( A => n40, B => n6, Z => neg_2a_12_port);
   U23 : XOR2_X1 port map( A => n44, B => n10, Z => neg_2a_16_port);
   U24 : XOR2_X1 port map( A => n47, B => n12, Z => neg_2a_19_port);
   U25 : XOR2_X1 port map( A => n37, B => n3, Z => neg_2a_9_port);
   U26 : XOR2_X1 port map( A => n39, B => n7, Z => neg_2a_11_port);
   U27 : XOR2_X1 port map( A => n43, B => n9, Z => neg_2a_15_port);
   U28 : XOR2_X1 port map( A => n46, B => n13, Z => neg_2a_18_port);
   U29 : XOR2_X1 port map( A => n38, B => n5, Z => neg_2a_10_port);
   U30 : XOR2_X1 port map( A => n42, B => n8, Z => neg_2a_14_port);
   U31 : XOR2_X1 port map( A => n45, B => n11, Z => neg_2a_17_port);
   U32 : XOR2_X1 port map( A => n49, B => n15, Z => neg_2a_21_port);
   U33 : XOR2_X1 port map( A => n41, B => n4, Z => neg_2a_13_port);
   U34 : XOR2_X1 port map( A => n48, B => n14, Z => neg_2a_20_port);
   U35 : INV_X1 port map( A => n33, ZN => pos_2a_22_port);
   U36 : INV_X1 port map( A => n33, ZN => pos_a_23_port);
   U37 : INV_X1 port map( A => a(14), ZN => n49);
   U38 : INV_X1 port map( A => a(13), ZN => n48);
   U39 : INV_X1 port map( A => a(12), ZN => n47);
   U40 : INV_X1 port map( A => a(11), ZN => n46);
   U41 : INV_X1 port map( A => a(10), ZN => n45);
   U42 : INV_X1 port map( A => a(9), ZN => n44);
   U43 : INV_X1 port map( A => a(8), ZN => n43);
   U44 : INV_X1 port map( A => a(7), ZN => n42);
   U45 : INV_X1 port map( A => a(6), ZN => n41);
   U46 : INV_X1 port map( A => a(5), ZN => n40);
   U47 : INV_X1 port map( A => a(4), ZN => n39);
   U48 : INV_X1 port map( A => a(3), ZN => n38);
   U49 : INV_X1 port map( A => a(2), ZN => n37);
   U50 : INV_X1 port map( A => a(1), ZN => n36);
   U51 : INV_X1 port map( A => a(0), ZN => n35);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT2 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT2;

architecture SYN_behavioral of shift_NBIT32_SHIFT2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_a_31, n1, neg_2a_20_port, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_6_port, neg_2a_10_port, 
      neg_2a_14_port, neg_2a_17_port, neg_2a_7_port, neg_2a_9_port, 
      neg_2a_13_port, neg_2a_16_port, neg_2a_8_port, neg_2a_12_port, 
      neg_2a_15_port, neg_2a_19_port, neg_2a_11_port, neg_2a_18_port, 
      pos_2a_20_port, pos_a_19_port, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49 : std_logic;

begin
   pos_a <= ( pos_a_19_port, pos_a_19_port, pos_a_19_port, pos_a_19_port, 
      pos_a_19_port, pos_a_19_port, pos_a_19_port, pos_a_19_port, pos_a_19_port
      , pos_a_19_port, pos_a_19_port, pos_a_19_port, pos_a_19_port, a(14), 
      a(13), a(12), a(11), a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), 
      a(2), a(1), a(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port );
   neg_a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_2a_20_port, neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, 
      neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, neg_2a_13_port, 
      neg_2a_12_port, neg_2a_11_port, neg_2a_10_port, neg_2a_9_port, 
      neg_2a_8_port, neg_2a_7_port, neg_2a_6_port, a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   pos_2a <= ( pos_2a_20_port, pos_2a_20_port, pos_2a_20_port, pos_2a_20_port, 
      pos_2a_20_port, pos_2a_20_port, pos_2a_20_port, pos_2a_20_port, 
      pos_2a_20_port, pos_2a_20_port, pos_2a_20_port, pos_2a_20_port, a(14), 
      a(13), a(12), a(11), a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), 
      a(2), a(1), a(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   neg_2a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_2a_20_port, 
      neg_2a_19_port, neg_2a_18_port, neg_2a_17_port, neg_2a_16_port, 
      neg_2a_15_port, neg_2a_14_port, neg_2a_13_port, neg_2a_12_port, 
      neg_2a_11_port, neg_2a_10_port, neg_2a_9_port, neg_2a_8_port, 
      neg_2a_7_port, neg_2a_6_port, a(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND2_X1 port map( A1 => n33, A2 => n16, ZN => n1);
   U3 : INV_X1 port map( A => n34, ZN => neg_a_31);
   U4 : XNOR2_X1 port map( A => n33, B => n1, ZN => n34);
   U5 : XOR2_X1 port map( A => n33, B => n16, Z => neg_2a_20_port);
   U6 : INV_X1 port map( A => a(15), ZN => n33);
   U7 : AND2_X1 port map( A1 => n36, A2 => n35, ZN => n3);
   U8 : AND2_X1 port map( A1 => n44, A2 => n11, ZN => n4);
   U9 : AND2_X1 port map( A1 => n37, A2 => n3, ZN => n5);
   U10 : AND2_X1 port map( A1 => n38, A2 => n5, ZN => n6);
   U11 : AND2_X1 port map( A1 => n39, A2 => n6, ZN => n7);
   U12 : AND2_X1 port map( A1 => n40, A2 => n7, ZN => n8);
   U13 : AND2_X1 port map( A1 => n41, A2 => n8, ZN => n9);
   U14 : AND2_X1 port map( A1 => n42, A2 => n9, ZN => n10);
   U15 : AND2_X1 port map( A1 => n43, A2 => n10, ZN => n11);
   U16 : AND2_X1 port map( A1 => n45, A2 => n4, ZN => n12);
   U17 : AND2_X1 port map( A1 => n46, A2 => n12, ZN => n13);
   U18 : AND2_X1 port map( A1 => n47, A2 => n13, ZN => n14);
   U19 : AND2_X1 port map( A1 => n48, A2 => n14, ZN => n15);
   U20 : AND2_X1 port map( A1 => n49, A2 => n15, ZN => n16);
   U21 : XOR2_X1 port map( A => n36, B => n35, Z => neg_2a_6_port);
   U22 : XOR2_X1 port map( A => n40, B => n7, Z => neg_2a_10_port);
   U23 : XOR2_X1 port map( A => n44, B => n11, Z => neg_2a_14_port);
   U24 : XOR2_X1 port map( A => n47, B => n13, Z => neg_2a_17_port);
   U25 : XOR2_X1 port map( A => n37, B => n3, Z => neg_2a_7_port);
   U26 : XOR2_X1 port map( A => n39, B => n6, Z => neg_2a_9_port);
   U27 : XOR2_X1 port map( A => n43, B => n10, Z => neg_2a_13_port);
   U28 : XOR2_X1 port map( A => n46, B => n12, Z => neg_2a_16_port);
   U29 : XOR2_X1 port map( A => n38, B => n5, Z => neg_2a_8_port);
   U30 : XOR2_X1 port map( A => n42, B => n9, Z => neg_2a_12_port);
   U31 : XOR2_X1 port map( A => n45, B => n4, Z => neg_2a_15_port);
   U32 : XOR2_X1 port map( A => n49, B => n15, Z => neg_2a_19_port);
   U33 : XOR2_X1 port map( A => n41, B => n8, Z => neg_2a_11_port);
   U34 : XOR2_X1 port map( A => n48, B => n14, Z => neg_2a_18_port);
   U35 : INV_X1 port map( A => n33, ZN => pos_2a_20_port);
   U36 : INV_X1 port map( A => n33, ZN => pos_a_19_port);
   U37 : INV_X1 port map( A => a(14), ZN => n49);
   U38 : INV_X1 port map( A => a(13), ZN => n48);
   U39 : INV_X1 port map( A => a(12), ZN => n47);
   U40 : INV_X1 port map( A => a(11), ZN => n46);
   U41 : INV_X1 port map( A => a(10), ZN => n45);
   U42 : INV_X1 port map( A => a(9), ZN => n44);
   U43 : INV_X1 port map( A => a(8), ZN => n43);
   U44 : INV_X1 port map( A => a(7), ZN => n42);
   U45 : INV_X1 port map( A => a(6), ZN => n41);
   U46 : INV_X1 port map( A => a(5), ZN => n40);
   U47 : INV_X1 port map( A => a(4), ZN => n39);
   U48 : INV_X1 port map( A => a(3), ZN => n38);
   U49 : INV_X1 port map( A => a(2), ZN => n37);
   U50 : INV_X1 port map( A => a(1), ZN => n36);
   U51 : INV_X1 port map( A => a(0), ZN => n35);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity rca_signed_NBIT32_0 is

   port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : out
         std_logic_vector (31 downto 0));

end rca_signed_NBIT32_0;

architecture SYN_Structural of rca_signed_NBIT32_0 is

   component fa_187
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_188
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_189
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_190
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_191
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_192
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_193
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_194
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_195
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_196
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_197
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_198
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_199
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_200
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_201
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_202
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_203
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_204
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_205
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_206
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_207
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_208
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_209
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_210
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_211
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_212
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_213
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_214
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_215
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_216
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component fa_0
      port( a, b, ci : in std_logic;  co, s : out std_logic);
   end component;
   
   component half_adder_0
      port( a, b : in std_logic;  co, s : out std_logic);
   end component;
   
   signal carry_s_30_port, carry_s_29_port, carry_s_28_port, carry_s_27_port, 
      carry_s_26_port, carry_s_25_port, carry_s_24_port, carry_s_23_port, 
      carry_s_22_port, carry_s_21_port, carry_s_20_port, carry_s_19_port, 
      carry_s_18_port, carry_s_17_port, carry_s_16_port, carry_s_15_port, 
      carry_s_14_port, carry_s_13_port, carry_s_12_port, carry_s_11_port, 
      carry_s_10_port, carry_s_9_port, carry_s_8_port, carry_s_7_port, 
      carry_s_6_port, carry_s_5_port, carry_s_4_port, carry_s_3_port, 
      carry_s_2_port, carry_s_1_port, carry_s_0_port : std_logic;

begin
   
   ha : half_adder_0 port map( a => a(0), b => b(0), co => carry_s_0_port, s =>
                           s(0));
   fa_i_1 : fa_0 port map( a => a(1), b => b(1), ci => carry_s_0_port, co => 
                           carry_s_1_port, s => s(1));
   fa_i_2 : fa_216 port map( a => a(2), b => b(2), ci => carry_s_1_port, co => 
                           carry_s_2_port, s => s(2));
   fa_i_3 : fa_215 port map( a => a(3), b => b(3), ci => carry_s_2_port, co => 
                           carry_s_3_port, s => s(3));
   fa_i_4 : fa_214 port map( a => a(4), b => b(4), ci => carry_s_3_port, co => 
                           carry_s_4_port, s => s(4));
   fa_i_5 : fa_213 port map( a => a(5), b => b(5), ci => carry_s_4_port, co => 
                           carry_s_5_port, s => s(5));
   fa_i_6 : fa_212 port map( a => a(6), b => b(6), ci => carry_s_5_port, co => 
                           carry_s_6_port, s => s(6));
   fa_i_7 : fa_211 port map( a => a(7), b => b(7), ci => carry_s_6_port, co => 
                           carry_s_7_port, s => s(7));
   fa_i_8 : fa_210 port map( a => a(8), b => b(8), ci => carry_s_7_port, co => 
                           carry_s_8_port, s => s(8));
   fa_i_9 : fa_209 port map( a => a(9), b => b(9), ci => carry_s_8_port, co => 
                           carry_s_9_port, s => s(9));
   fa_i_10 : fa_208 port map( a => a(10), b => b(10), ci => carry_s_9_port, co 
                           => carry_s_10_port, s => s(10));
   fa_i_11 : fa_207 port map( a => a(11), b => b(11), ci => carry_s_10_port, co
                           => carry_s_11_port, s => s(11));
   fa_i_12 : fa_206 port map( a => a(12), b => b(12), ci => carry_s_11_port, co
                           => carry_s_12_port, s => s(12));
   fa_i_13 : fa_205 port map( a => a(13), b => b(13), ci => carry_s_12_port, co
                           => carry_s_13_port, s => s(13));
   fa_i_14 : fa_204 port map( a => a(14), b => b(14), ci => carry_s_13_port, co
                           => carry_s_14_port, s => s(14));
   fa_i_15 : fa_203 port map( a => a(15), b => b(15), ci => carry_s_14_port, co
                           => carry_s_15_port, s => s(15));
   fa_i_16 : fa_202 port map( a => a(16), b => b(16), ci => carry_s_15_port, co
                           => carry_s_16_port, s => s(16));
   fa_i_17 : fa_201 port map( a => a(17), b => b(17), ci => carry_s_16_port, co
                           => carry_s_17_port, s => s(17));
   fa_i_18 : fa_200 port map( a => a(18), b => b(18), ci => carry_s_17_port, co
                           => carry_s_18_port, s => s(18));
   fa_i_19 : fa_199 port map( a => a(19), b => b(19), ci => carry_s_18_port, co
                           => carry_s_19_port, s => s(19));
   fa_i_20 : fa_198 port map( a => a(20), b => b(20), ci => carry_s_19_port, co
                           => carry_s_20_port, s => s(20));
   fa_i_21 : fa_197 port map( a => a(21), b => b(21), ci => carry_s_20_port, co
                           => carry_s_21_port, s => s(21));
   fa_i_22 : fa_196 port map( a => a(22), b => b(22), ci => carry_s_21_port, co
                           => carry_s_22_port, s => s(22));
   fa_i_23 : fa_195 port map( a => a(23), b => b(23), ci => carry_s_22_port, co
                           => carry_s_23_port, s => s(23));
   fa_i_24 : fa_194 port map( a => a(24), b => b(24), ci => carry_s_23_port, co
                           => carry_s_24_port, s => s(24));
   fa_i_25 : fa_193 port map( a => a(25), b => b(25), ci => carry_s_24_port, co
                           => carry_s_25_port, s => s(25));
   fa_i_26 : fa_192 port map( a => a(26), b => b(26), ci => carry_s_25_port, co
                           => carry_s_26_port, s => s(26));
   fa_i_27 : fa_191 port map( a => a(27), b => b(27), ci => carry_s_26_port, co
                           => carry_s_27_port, s => s(27));
   fa_i_28 : fa_190 port map( a => a(28), b => b(28), ci => carry_s_27_port, co
                           => carry_s_28_port, s => s(28));
   fa_i_29 : fa_189 port map( a => a(29), b => b(29), ci => carry_s_28_port, co
                           => carry_s_29_port, s => s(29));
   fa_i_30 : fa_188 port map( a => a(30), b => b(30), ci => carry_s_29_port, co
                           => carry_s_30_port, s => s(30));
   fa_i_31 : fa_187 port map( a => a(31), b => b(31), ci => carry_s_30_port, co
                           => c, s => s(31));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT1 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT1;

architecture SYN_behavioral of shift_NBIT32_SHIFT1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_a_31, n1, neg_2a_18_port, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_4_port, neg_2a_8_port, 
      neg_2a_12_port, neg_2a_15_port, neg_2a_5_port, neg_2a_7_port, 
      neg_2a_11_port, neg_2a_14_port, neg_2a_6_port, neg_2a_10_port, 
      neg_2a_13_port, neg_2a_17_port, neg_2a_9_port, neg_2a_16_port, 
      pos_2a_18_port, pos_2a_30_port, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49 : std_logic;

begin
   pos_a <= ( pos_2a_30_port, pos_2a_18_port, pos_2a_30_port, pos_2a_18_port, 
      pos_2a_30_port, pos_2a_30_port, pos_2a_30_port, pos_2a_30_port, 
      pos_2a_30_port, pos_2a_30_port, pos_2a_30_port, pos_2a_30_port, 
      pos_2a_30_port, pos_2a_30_port, pos_2a_30_port, a(14), a(13), a(12), 
      a(11), a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0),
      X_Logic0_port, X_Logic0_port );
   neg_a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_2a_18_port, neg_2a_17_port, neg_2a_16_port, neg_2a_15_port,
      neg_2a_14_port, neg_2a_13_port, neg_2a_12_port, neg_2a_11_port, 
      neg_2a_10_port, neg_2a_9_port, neg_2a_8_port, neg_2a_7_port, 
      neg_2a_6_port, neg_2a_5_port, neg_2a_4_port, a(0), X_Logic0_port, 
      X_Logic0_port );
   pos_2a <= ( pos_2a_30_port, pos_2a_30_port, pos_2a_18_port, pos_2a_18_port, 
      pos_2a_18_port, pos_2a_18_port, pos_2a_18_port, pos_2a_18_port, 
      pos_2a_18_port, pos_2a_18_port, pos_2a_18_port, pos_2a_18_port, 
      pos_2a_18_port, pos_2a_18_port, a(14), a(13), a(12), a(11), a(10), a(9), 
      a(8), a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   neg_2a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_2a_18_port, neg_2a_17_port, neg_2a_16_port, neg_2a_15_port, 
      neg_2a_14_port, neg_2a_13_port, neg_2a_12_port, neg_2a_11_port, 
      neg_2a_10_port, neg_2a_9_port, neg_2a_8_port, neg_2a_7_port, 
      neg_2a_6_port, neg_2a_5_port, neg_2a_4_port, a(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND2_X1 port map( A1 => n33, A2 => n16, ZN => n1);
   U3 : XNOR2_X1 port map( A => n33, B => n1, ZN => n34);
   U4 : XOR2_X1 port map( A => n33, B => n16, Z => neg_2a_18_port);
   U5 : INV_X1 port map( A => a(15), ZN => n33);
   U6 : AND2_X1 port map( A1 => n36, A2 => n35, ZN => n3);
   U7 : AND2_X1 port map( A1 => n37, A2 => n3, ZN => n4);
   U8 : AND2_X1 port map( A1 => n38, A2 => n4, ZN => n5);
   U9 : AND2_X1 port map( A1 => n40, A2 => n7, ZN => n6);
   U10 : AND2_X1 port map( A1 => n39, A2 => n5, ZN => n7);
   U11 : AND2_X1 port map( A1 => n42, A2 => n15, ZN => n8);
   U12 : AND2_X1 port map( A1 => n43, A2 => n8, ZN => n9);
   U13 : AND2_X1 port map( A1 => n44, A2 => n9, ZN => n10);
   U14 : AND2_X1 port map( A1 => n47, A2 => n13, ZN => n11);
   U15 : AND2_X1 port map( A1 => n45, A2 => n10, ZN => n12);
   U16 : AND2_X1 port map( A1 => n46, A2 => n12, ZN => n13);
   U17 : AND2_X1 port map( A1 => n48, A2 => n11, ZN => n14);
   U18 : AND2_X1 port map( A1 => n41, A2 => n6, ZN => n15);
   U19 : AND2_X1 port map( A1 => n49, A2 => n14, ZN => n16);
   U20 : XOR2_X1 port map( A => n36, B => n35, Z => neg_2a_4_port);
   U21 : XOR2_X1 port map( A => n40, B => n7, Z => neg_2a_8_port);
   U22 : XOR2_X1 port map( A => n44, B => n9, Z => neg_2a_12_port);
   U23 : XOR2_X1 port map( A => n47, B => n13, Z => neg_2a_15_port);
   U24 : XOR2_X1 port map( A => n37, B => n3, Z => neg_2a_5_port);
   U25 : XOR2_X1 port map( A => n39, B => n5, Z => neg_2a_7_port);
   U26 : XOR2_X1 port map( A => n43, B => n8, Z => neg_2a_11_port);
   U27 : XOR2_X1 port map( A => n46, B => n12, Z => neg_2a_14_port);
   U28 : XOR2_X1 port map( A => n38, B => n4, Z => neg_2a_6_port);
   U29 : XOR2_X1 port map( A => n42, B => n15, Z => neg_2a_10_port);
   U30 : XOR2_X1 port map( A => n45, B => n10, Z => neg_2a_13_port);
   U31 : XOR2_X1 port map( A => n49, B => n14, Z => neg_2a_17_port);
   U32 : XOR2_X1 port map( A => n41, B => n6, Z => neg_2a_9_port);
   U33 : XOR2_X1 port map( A => n48, B => n11, Z => neg_2a_16_port);
   U34 : INV_X1 port map( A => n33, ZN => pos_2a_18_port);
   U35 : INV_X1 port map( A => n33, ZN => pos_2a_30_port);
   U36 : INV_X2 port map( A => n34, ZN => neg_a_31);
   U37 : INV_X1 port map( A => a(14), ZN => n49);
   U38 : INV_X1 port map( A => a(13), ZN => n48);
   U39 : INV_X1 port map( A => a(12), ZN => n47);
   U40 : INV_X1 port map( A => a(11), ZN => n46);
   U41 : INV_X1 port map( A => a(10), ZN => n45);
   U42 : INV_X1 port map( A => a(9), ZN => n44);
   U43 : INV_X1 port map( A => a(8), ZN => n43);
   U44 : INV_X1 port map( A => a(7), ZN => n42);
   U45 : INV_X1 port map( A => a(6), ZN => n41);
   U46 : INV_X1 port map( A => a(5), ZN => n40);
   U47 : INV_X1 port map( A => a(4), ZN => n39);
   U48 : INV_X1 port map( A => a(3), ZN => n38);
   U49 : INV_X1 port map( A => a(2), ZN => n37);
   U50 : INV_X1 port map( A => a(1), ZN => n36);
   U51 : INV_X1 port map( A => a(0), ZN => n35);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity vp_NBIT32_0 is

   port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  sel
         : in std_logic_vector (2 downto 0);  s_out : out std_logic_vector (31 
         downto 0));

end vp_NBIT32_0;

architecture SYN_behavioral of vp_NBIT32_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n70, A2 => n71, ZN => n5);
   U3 : AND3_X2 port map( A1 => sel(1), A2 => n71, A3 => sel(0), ZN => n7);
   U4 : AND2_X2 port map( A1 => sel(2), A2 => n70, ZN => n6);
   U5 : OR3_X1 port map( A1 => sel(0), A2 => sel(1), A3 => n71, ZN => n4);
   U6 : INV_X2 port map( A => n4, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => s_out(9));
   U8 : AOI22_X1 port map( A1 => neg_2a(9), A2 => n1, B1 => pos_a(9), B2 => n5,
                           ZN => n3);
   U9 : AOI22_X1 port map( A1 => neg_a(9), A2 => n6, B1 => pos_2a(9), B2 => n7,
                           ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => s_out(8));
   U11 : AOI22_X1 port map( A1 => neg_2a(8), A2 => n1, B1 => pos_a(8), B2 => n5
                           , ZN => n9);
   U12 : AOI22_X1 port map( A1 => neg_a(8), A2 => n6, B1 => pos_2a(8), B2 => n7
                           , ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => s_out(7));
   U14 : AOI22_X1 port map( A1 => neg_2a(7), A2 => n1, B1 => pos_a(7), B2 => n5
                           , ZN => n11);
   U15 : AOI22_X1 port map( A1 => neg_a(7), A2 => n6, B1 => pos_2a(7), B2 => n7
                           , ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => s_out(6));
   U17 : AOI22_X1 port map( A1 => neg_2a(6), A2 => n1, B1 => pos_a(6), B2 => n5
                           , ZN => n13);
   U18 : AOI22_X1 port map( A1 => neg_a(6), A2 => n6, B1 => pos_2a(6), B2 => n7
                           , ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => s_out(5));
   U20 : AOI22_X1 port map( A1 => neg_2a(5), A2 => n1, B1 => pos_a(5), B2 => n5
                           , ZN => n15);
   U21 : AOI22_X1 port map( A1 => neg_a(5), A2 => n6, B1 => pos_2a(5), B2 => n7
                           , ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => s_out(4));
   U23 : AOI22_X1 port map( A1 => neg_2a(4), A2 => n1, B1 => pos_a(4), B2 => n5
                           , ZN => n17);
   U24 : AOI22_X1 port map( A1 => neg_a(4), A2 => n6, B1 => pos_2a(4), B2 => n7
                           , ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => s_out(3));
   U26 : AOI22_X1 port map( A1 => neg_2a(3), A2 => n1, B1 => pos_a(3), B2 => n5
                           , ZN => n19);
   U27 : AOI22_X1 port map( A1 => neg_a(3), A2 => n6, B1 => pos_2a(3), B2 => n7
                           , ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => s_out(31));
   U29 : AOI22_X1 port map( A1 => neg_2a(31), A2 => n1, B1 => pos_a(31), B2 => 
                           n5, ZN => n21);
   U30 : AOI22_X1 port map( A1 => neg_a(31), A2 => n6, B1 => pos_2a(31), B2 => 
                           n7, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => s_out(30));
   U32 : AOI22_X1 port map( A1 => neg_2a(30), A2 => n1, B1 => pos_a(30), B2 => 
                           n5, ZN => n23);
   U33 : AOI22_X1 port map( A1 => neg_a(30), A2 => n6, B1 => pos_2a(30), B2 => 
                           n7, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => s_out(2));
   U35 : AOI22_X1 port map( A1 => neg_2a(2), A2 => n1, B1 => pos_a(2), B2 => n5
                           , ZN => n25);
   U36 : AOI22_X1 port map( A1 => neg_a(2), A2 => n6, B1 => pos_2a(2), B2 => n7
                           , ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => s_out(29));
   U38 : AOI22_X1 port map( A1 => neg_2a(29), A2 => n1, B1 => pos_a(29), B2 => 
                           n5, ZN => n27);
   U39 : AOI22_X1 port map( A1 => neg_a(29), A2 => n6, B1 => pos_2a(29), B2 => 
                           n7, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => s_out(28));
   U41 : AOI22_X1 port map( A1 => neg_2a(28), A2 => n1, B1 => pos_a(28), B2 => 
                           n5, ZN => n29);
   U42 : AOI22_X1 port map( A1 => neg_a(28), A2 => n6, B1 => pos_2a(28), B2 => 
                           n7, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => s_out(27));
   U44 : AOI22_X1 port map( A1 => neg_2a(27), A2 => n1, B1 => pos_a(27), B2 => 
                           n5, ZN => n31);
   U45 : AOI22_X1 port map( A1 => neg_a(27), A2 => n6, B1 => pos_2a(27), B2 => 
                           n7, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => s_out(26));
   U47 : AOI22_X1 port map( A1 => neg_2a(26), A2 => n1, B1 => pos_a(26), B2 => 
                           n5, ZN => n33);
   U48 : AOI22_X1 port map( A1 => neg_a(26), A2 => n6, B1 => pos_2a(26), B2 => 
                           n7, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => s_out(25));
   U50 : AOI22_X1 port map( A1 => neg_2a(25), A2 => n1, B1 => pos_a(25), B2 => 
                           n5, ZN => n35);
   U51 : AOI22_X1 port map( A1 => neg_a(25), A2 => n6, B1 => pos_2a(25), B2 => 
                           n7, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => s_out(24));
   U53 : AOI22_X1 port map( A1 => neg_2a(24), A2 => n1, B1 => pos_a(24), B2 => 
                           n5, ZN => n37);
   U54 : AOI22_X1 port map( A1 => neg_a(24), A2 => n6, B1 => pos_2a(24), B2 => 
                           n7, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => s_out(23));
   U56 : AOI22_X1 port map( A1 => neg_2a(23), A2 => n1, B1 => pos_a(23), B2 => 
                           n5, ZN => n39);
   U57 : AOI22_X1 port map( A1 => neg_a(23), A2 => n6, B1 => pos_2a(23), B2 => 
                           n7, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => s_out(22));
   U59 : AOI22_X1 port map( A1 => neg_2a(22), A2 => n1, B1 => pos_a(22), B2 => 
                           n5, ZN => n41);
   U60 : AOI22_X1 port map( A1 => neg_a(22), A2 => n6, B1 => pos_2a(22), B2 => 
                           n7, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => s_out(21));
   U62 : AOI22_X1 port map( A1 => neg_2a(21), A2 => n1, B1 => pos_a(21), B2 => 
                           n5, ZN => n43);
   U63 : AOI22_X1 port map( A1 => neg_a(21), A2 => n6, B1 => pos_2a(21), B2 => 
                           n7, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => s_out(20));
   U65 : AOI22_X1 port map( A1 => neg_2a(20), A2 => n1, B1 => pos_a(20), B2 => 
                           n5, ZN => n45);
   U66 : AOI22_X1 port map( A1 => neg_a(20), A2 => n6, B1 => pos_2a(20), B2 => 
                           n7, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => s_out(1));
   U68 : AOI22_X1 port map( A1 => neg_2a(1), A2 => n1, B1 => pos_a(1), B2 => n5
                           , ZN => n47);
   U69 : AOI22_X1 port map( A1 => neg_a(1), A2 => n6, B1 => pos_2a(1), B2 => n7
                           , ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => s_out(19));
   U71 : AOI22_X1 port map( A1 => neg_2a(19), A2 => n1, B1 => pos_a(19), B2 => 
                           n5, ZN => n49);
   U72 : AOI22_X1 port map( A1 => neg_a(19), A2 => n6, B1 => pos_2a(19), B2 => 
                           n7, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => s_out(18));
   U74 : AOI22_X1 port map( A1 => neg_2a(18), A2 => n1, B1 => pos_a(18), B2 => 
                           n5, ZN => n51);
   U75 : AOI22_X1 port map( A1 => neg_a(18), A2 => n6, B1 => pos_2a(18), B2 => 
                           n7, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => s_out(17));
   U77 : AOI22_X1 port map( A1 => neg_2a(17), A2 => n1, B1 => pos_a(17), B2 => 
                           n5, ZN => n53);
   U78 : AOI22_X1 port map( A1 => neg_a(17), A2 => n6, B1 => pos_2a(17), B2 => 
                           n7, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => s_out(16));
   U80 : AOI22_X1 port map( A1 => neg_2a(16), A2 => n1, B1 => pos_a(16), B2 => 
                           n5, ZN => n55);
   U81 : AOI22_X1 port map( A1 => neg_a(16), A2 => n6, B1 => pos_2a(16), B2 => 
                           n7, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => s_out(15));
   U83 : AOI22_X1 port map( A1 => neg_2a(15), A2 => n1, B1 => pos_a(15), B2 => 
                           n5, ZN => n57);
   U84 : AOI22_X1 port map( A1 => neg_a(15), A2 => n6, B1 => pos_2a(15), B2 => 
                           n7, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => s_out(14));
   U86 : AOI22_X1 port map( A1 => neg_2a(14), A2 => n1, B1 => pos_a(14), B2 => 
                           n5, ZN => n59);
   U87 : AOI22_X1 port map( A1 => neg_a(14), A2 => n6, B1 => pos_2a(14), B2 => 
                           n7, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => s_out(13));
   U89 : AOI22_X1 port map( A1 => neg_2a(13), A2 => n1, B1 => pos_a(13), B2 => 
                           n5, ZN => n61);
   U90 : AOI22_X1 port map( A1 => neg_a(13), A2 => n6, B1 => pos_2a(13), B2 => 
                           n7, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => s_out(12));
   U92 : AOI22_X1 port map( A1 => neg_2a(12), A2 => n1, B1 => pos_a(12), B2 => 
                           n5, ZN => n63);
   U93 : AOI22_X1 port map( A1 => neg_a(12), A2 => n6, B1 => pos_2a(12), B2 => 
                           n7, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => s_out(11));
   U95 : AOI22_X1 port map( A1 => neg_2a(11), A2 => n1, B1 => pos_a(11), B2 => 
                           n5, ZN => n65);
   U96 : AOI22_X1 port map( A1 => neg_a(11), A2 => n6, B1 => pos_2a(11), B2 => 
                           n7, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => s_out(10));
   U98 : AOI22_X1 port map( A1 => neg_2a(10), A2 => n1, B1 => pos_a(10), B2 => 
                           n5, ZN => n67);
   U99 : AOI22_X1 port map( A1 => neg_a(10), A2 => n6, B1 => pos_2a(10), B2 => 
                           n7, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => s_out(0));
   U101 : AOI22_X1 port map( A1 => neg_2a(0), A2 => n1, B1 => pos_a(0), B2 => 
                           n5, ZN => n69);
   U102 : AOI22_X1 port map( A1 => neg_a(0), A2 => n6, B1 => pos_2a(0), B2 => 
                           n7, ZN => n68);
   U103 : INV_X1 port map( A => sel(2), ZN => n71);
   U104 : XOR2_X1 port map( A => sel(0), B => sel(1), Z => n70);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shift_NBIT32_SHIFT0 is

   port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, neg_2a :
         out std_logic_vector (31 downto 0));

end shift_NBIT32_SHIFT0;

architecture SYN_behavioral of shift_NBIT32_SHIFT0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, neg_a_31, n1, neg_2a_16_port, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, neg_2a_2_port, neg_2a_6_port, 
      neg_2a_10_port, neg_2a_13_port, neg_2a_3_port, neg_2a_5_port, 
      neg_2a_9_port, neg_2a_12_port, neg_2a_4_port, neg_2a_8_port, 
      neg_2a_11_port, neg_2a_15_port, neg_2a_7_port, neg_2a_14_port, 
      pos_2a_16_port, pos_2a_28_port, pos_a_23_port, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50 : std_logic;

begin
   pos_a <= ( pos_a_23_port, pos_a_23_port, pos_a_23_port, pos_a_23_port, 
      pos_a_23_port, pos_a_23_port, pos_a_23_port, pos_a_23_port, pos_a_23_port
      , pos_2a_28_port, pos_2a_28_port, pos_2a_28_port, pos_2a_28_port, 
      pos_2a_28_port, pos_2a_28_port, pos_2a_28_port, pos_2a_28_port, a(14), 
      a(13), a(12), a(11), a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), 
      a(2), a(1), a(0) );
   neg_a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_2a_16_port, neg_2a_15_port, 
      neg_2a_14_port, neg_2a_13_port, neg_2a_12_port, neg_2a_11_port, 
      neg_2a_10_port, neg_2a_9_port, neg_2a_8_port, neg_2a_7_port, 
      neg_2a_6_port, neg_2a_5_port, neg_2a_4_port, neg_2a_3_port, neg_2a_2_port
      , a(0) );
   pos_2a <= ( pos_2a_28_port, pos_2a_28_port, pos_2a_28_port, pos_2a_28_port, 
      pos_2a_16_port, pos_2a_16_port, pos_2a_16_port, pos_2a_16_port, 
      pos_2a_16_port, pos_2a_16_port, pos_2a_16_port, pos_2a_16_port, 
      pos_2a_16_port, pos_2a_16_port, pos_2a_16_port, pos_2a_16_port, a(14), 
      a(13), a(12), a(11), a(10), a(9), a(8), a(7), a(6), a(5), a(4), a(3), 
      a(2), a(1), a(0), X_Logic0_port );
   neg_2a <= ( neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, neg_a_31, 
      neg_a_31, neg_a_31, neg_2a_16_port, neg_2a_15_port, neg_2a_14_port, 
      neg_2a_13_port, neg_2a_12_port, neg_2a_11_port, neg_2a_10_port, 
      neg_2a_9_port, neg_2a_8_port, neg_2a_7_port, neg_2a_6_port, neg_2a_5_port
      , neg_2a_4_port, neg_2a_3_port, neg_2a_2_port, a(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND2_X1 port map( A1 => n34, A2 => n16, ZN => n1);
   U3 : XNOR2_X1 port map( A => n34, B => n1, ZN => n35);
   U4 : XOR2_X1 port map( A => n34, B => n16, Z => neg_2a_16_port);
   U5 : INV_X1 port map( A => a(15), ZN => n34);
   U6 : AND2_X1 port map( A1 => n37, A2 => n36, ZN => n3);
   U7 : AND2_X1 port map( A1 => n38, A2 => n3, ZN => n4);
   U8 : AND2_X1 port map( A1 => n39, A2 => n4, ZN => n5);
   U9 : AND2_X1 port map( A1 => n40, A2 => n5, ZN => n6);
   U10 : AND2_X1 port map( A1 => n41, A2 => n6, ZN => n7);
   U11 : AND2_X1 port map( A1 => n48, A2 => n14, ZN => n8);
   U12 : AND2_X1 port map( A1 => n42, A2 => n7, ZN => n9);
   U13 : AND2_X1 port map( A1 => n43, A2 => n9, ZN => n10);
   U14 : AND2_X1 port map( A1 => n44, A2 => n10, ZN => n11);
   U15 : AND2_X1 port map( A1 => n45, A2 => n11, ZN => n12);
   U16 : AND2_X1 port map( A1 => n46, A2 => n12, ZN => n13);
   U17 : AND2_X1 port map( A1 => n47, A2 => n13, ZN => n14);
   U18 : AND2_X1 port map( A1 => n49, A2 => n8, ZN => n15);
   U19 : AND2_X1 port map( A1 => n50, A2 => n15, ZN => n16);
   U20 : XOR2_X1 port map( A => n37, B => n36, Z => neg_2a_2_port);
   U21 : XOR2_X1 port map( A => n41, B => n6, Z => neg_2a_6_port);
   U22 : XOR2_X1 port map( A => n45, B => n11, Z => neg_2a_10_port);
   U23 : XOR2_X1 port map( A => n48, B => n14, Z => neg_2a_13_port);
   U24 : XOR2_X1 port map( A => n38, B => n3, Z => neg_2a_3_port);
   U25 : XOR2_X1 port map( A => n40, B => n5, Z => neg_2a_5_port);
   U26 : XOR2_X1 port map( A => n44, B => n10, Z => neg_2a_9_port);
   U27 : XOR2_X1 port map( A => n47, B => n13, Z => neg_2a_12_port);
   U28 : XOR2_X1 port map( A => n39, B => n4, Z => neg_2a_4_port);
   U29 : XOR2_X1 port map( A => n43, B => n9, Z => neg_2a_8_port);
   U30 : XOR2_X1 port map( A => n46, B => n12, Z => neg_2a_11_port);
   U31 : XOR2_X1 port map( A => n50, B => n15, Z => neg_2a_15_port);
   U32 : XOR2_X1 port map( A => n42, B => n7, Z => neg_2a_7_port);
   U33 : XOR2_X1 port map( A => n49, B => n8, Z => neg_2a_14_port);
   U34 : INV_X1 port map( A => n34, ZN => pos_2a_16_port);
   U35 : INV_X1 port map( A => n34, ZN => pos_2a_28_port);
   U36 : INV_X1 port map( A => n34, ZN => pos_a_23_port);
   U37 : INV_X2 port map( A => n35, ZN => neg_a_31);
   U38 : INV_X1 port map( A => a(14), ZN => n50);
   U39 : INV_X1 port map( A => a(13), ZN => n49);
   U40 : INV_X1 port map( A => a(12), ZN => n48);
   U41 : INV_X1 port map( A => a(11), ZN => n47);
   U42 : INV_X1 port map( A => a(10), ZN => n46);
   U43 : INV_X1 port map( A => a(9), ZN => n45);
   U44 : INV_X1 port map( A => a(8), ZN => n44);
   U45 : INV_X1 port map( A => a(7), ZN => n43);
   U46 : INV_X1 port map( A => a(6), ZN => n42);
   U47 : INV_X1 port map( A => a(5), ZN => n41);
   U48 : INV_X1 port map( A => a(4), ZN => n40);
   U49 : INV_X1 port map( A => a(3), ZN => n39);
   U50 : INV_X1 port map( A => a(2), ZN => n38);
   U51 : INV_X1 port map( A => a(1), ZN => n37);
   U52 : INV_X1 port map( A => a(0), ZN => n36);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity carry_select_adder_n_bit4_0 is

   port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (3 downto 0);  carry_out, 
         overflow : out std_logic);

end carry_select_adder_n_bit4_0;

architecture SYN_specification of carry_select_adder_n_bit4_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_15
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component ripple_carry_adder_n_bit4_0
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ovf_1_port, ovf_0_port, cout_1_port, 
      cout_0_port, sumsig_7_port, sumsig_6_port, sumsig_5_port, sumsig_4_port, 
      sumsig_3_port, sumsig_2_port, sumsig_1_port, sumsig_0_port : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_0 : ripple_carry_adder_n_bit4_0 port map( operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic0_port, sum(3) => sumsig_3_port, sum(2) => 
                           sumsig_2_port, sum(1) => sumsig_1_port, sum(0) => 
                           sumsig_0_port, carry_out => cout_0_port, overflow =>
                           ovf_0_port);
   rca_1 : ripple_carry_adder_n_bit4_15 port map( operand_1(3) => operand_1(3),
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => 
                           X_Logic1_port, sum(3) => sumsig_7_port, sum(2) => 
                           sumsig_6_port, sum(1) => sumsig_5_port, sum(0) => 
                           sumsig_4_port, carry_out => cout_1_port, overflow =>
                           ovf_1_port);
   U3 : MUX2_X1 port map( A => cout_0_port, B => cout_1_port, S => carry_in, Z 
                           => carry_out);
   U4 : MUX2_X1 port map( A => ovf_0_port, B => ovf_1_port, S => carry_in, Z =>
                           overflow);
   U5 : MUX2_X1 port map( A => sumsig_3_port, B => sumsig_7_port, S => carry_in
                           , Z => sum(3));
   U6 : MUX2_X1 port map( A => sumsig_2_port, B => sumsig_6_port, S => carry_in
                           , Z => sum(2));
   U7 : MUX2_X1 port map( A => sumsig_1_port, B => sumsig_5_port, S => carry_in
                           , Z => sum(1));
   U8 : MUX2_X1 port map( A => sumsig_0_port, B => sumsig_4_port, S => carry_in
                           , Z => sum(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity sparse_tree_carry_generator_n_bit32 is

   port( operand_1, operand_2 : in std_logic_vector (31 downto 0);  carry_in : 
         in std_logic;  carry_out : out std_logic_vector (7 downto 0));

end sparse_tree_carry_generator_n_bit32;

architecture SYN_specification of sparse_tree_carry_generator_n_bit32 is

   component g_block_1
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component g_block_2
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component g_block_3
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component g_block_4
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component pg_block_1
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_2
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component g_block_5
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component g_block_6
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component pg_block_3
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_4
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_5
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component g_block_7
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component pg_block_6
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_7
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_8
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_9
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_10
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_11
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_12
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component g_block_0
      port( Gik, Pik, Gk1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component pg_block_13
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_14
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_15
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_16
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_17
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_18
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_19
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_20
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_21
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_22
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_23
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_24
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_25
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_26
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component pg_block_0
      port( Gik, Pik, Gk1j, Pk1j : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component g_block_carry
      port( Gik, Pik, Gk1j, Pk1j, carry_in : in std_logic;  Gij : out std_logic
            );
   end component;
   
   component pg_network_n_bit32
      port( operand_1, operand_2 : in std_logic_vector (32 downto 1);  p, g : 
            out std_logic_vector (32 downto 1));
   end component;
   
   signal carry_out_7_port, carry_out_6_port, carry_out_5_port, 
      carry_out_4_port, carry_out_3_port, carry_out_2_port, carry_out_1_port, 
      carry_out_0_port, p_31_port, p_30_port, p_29_port, p_28_port, p_27_port, 
      p_26_port, p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, 
      p_20_port, p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, 
      p_14_port, p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port
      , p_7_port, p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, 
      p_0_port, g_31_port, g_30_port, g_29_port, g_28_port, g_27_port, 
      g_26_port, g_25_port, g_24_port, g_23_port, g_22_port, g_21_port, 
      g_20_port, g_19_port, g_18_port, g_17_port, g_16_port, g_15_port, 
      g_14_port, g_13_port, g_12_port, g_11_port, g_10_port, g_9_port, g_8_port
      , g_7_port, g_6_port, g_5_port, g_4_port, g_3_port, g_2_port, g_1_port, 
      g_0_port, g_matrix_0_15_port, g_matrix_0_14_port, g_matrix_0_13_port, 
      g_matrix_0_12_port, g_matrix_0_11_port, g_matrix_0_10_port, 
      g_matrix_0_9_port, g_matrix_0_8_port, g_matrix_0_7_port, 
      g_matrix_0_6_port, g_matrix_0_5_port, g_matrix_0_4_port, 
      g_matrix_0_3_port, g_matrix_0_2_port, g_matrix_0_1_port, 
      g_matrix_0_0_port, g_matrix_1_7_port, g_matrix_1_6_port, 
      g_matrix_1_5_port, g_matrix_1_4_port, g_matrix_1_3_port, 
      g_matrix_1_2_port, g_matrix_1_1_port, g_matrix_2_7_port, 
      g_matrix_2_5_port, g_matrix_2_3_port, g_matrix_3_7_port, 
      g_matrix_3_6_port, p_matrix_0_15_port, p_matrix_0_14_port, 
      p_matrix_0_13_port, p_matrix_0_12_port, p_matrix_0_11_port, 
      p_matrix_0_10_port, p_matrix_0_9_port, p_matrix_0_8_port, 
      p_matrix_0_7_port, p_matrix_0_6_port, p_matrix_0_5_port, 
      p_matrix_0_4_port, p_matrix_0_3_port, p_matrix_0_2_port, 
      p_matrix_0_1_port, p_matrix_1_7_port, p_matrix_1_6_port, 
      p_matrix_1_5_port, p_matrix_1_4_port, p_matrix_1_3_port, 
      p_matrix_1_2_port, p_matrix_1_1_port, p_matrix_2_7_port, 
      p_matrix_2_5_port, p_matrix_2_3_port, p_matrix_3_7_port, 
      p_matrix_3_6_port : std_logic;

begin
   carry_out <= ( carry_out_7_port, carry_out_6_port, carry_out_5_port, 
      carry_out_4_port, carry_out_3_port, carry_out_2_port, carry_out_1_port, 
      carry_out_0_port );
   
   pgnetwork : pg_network_n_bit32 port map( operand_1(32) => operand_1(31), 
                           operand_1(31) => operand_1(30), operand_1(30) => 
                           operand_1(29), operand_1(29) => operand_1(28), 
                           operand_1(28) => operand_1(27), operand_1(27) => 
                           operand_1(26), operand_1(26) => operand_1(25), 
                           operand_1(25) => operand_1(24), operand_1(24) => 
                           operand_1(23), operand_1(23) => operand_1(22), 
                           operand_1(22) => operand_1(21), operand_1(21) => 
                           operand_1(20), operand_1(20) => operand_1(19), 
                           operand_1(19) => operand_1(18), operand_1(18) => 
                           operand_1(17), operand_1(17) => operand_1(16), 
                           operand_1(16) => operand_1(15), operand_1(15) => 
                           operand_1(14), operand_1(14) => operand_1(13), 
                           operand_1(13) => operand_1(12), operand_1(12) => 
                           operand_1(11), operand_1(11) => operand_1(10), 
                           operand_1(10) => operand_1(9), operand_1(9) => 
                           operand_1(8), operand_1(8) => operand_1(7), 
                           operand_1(7) => operand_1(6), operand_1(6) => 
                           operand_1(5), operand_1(5) => operand_1(4), 
                           operand_1(4) => operand_1(3), operand_1(3) => 
                           operand_1(2), operand_1(2) => operand_1(1), 
                           operand_1(1) => operand_1(0), operand_2(32) => 
                           operand_2(31), operand_2(31) => operand_2(30), 
                           operand_2(30) => operand_2(29), operand_2(29) => 
                           operand_2(28), operand_2(28) => operand_2(27), 
                           operand_2(27) => operand_2(26), operand_2(26) => 
                           operand_2(25), operand_2(25) => operand_2(24), 
                           operand_2(24) => operand_2(23), operand_2(23) => 
                           operand_2(22), operand_2(22) => operand_2(21), 
                           operand_2(21) => operand_2(20), operand_2(20) => 
                           operand_2(19), operand_2(19) => operand_2(18), 
                           operand_2(18) => operand_2(17), operand_2(17) => 
                           operand_2(16), operand_2(16) => operand_2(15), 
                           operand_2(15) => operand_2(14), operand_2(14) => 
                           operand_2(13), operand_2(13) => operand_2(12), 
                           operand_2(12) => operand_2(11), operand_2(11) => 
                           operand_2(10), operand_2(10) => operand_2(9), 
                           operand_2(9) => operand_2(8), operand_2(8) => 
                           operand_2(7), operand_2(7) => operand_2(6), 
                           operand_2(6) => operand_2(5), operand_2(5) => 
                           operand_2(4), operand_2(4) => operand_2(3), 
                           operand_2(3) => operand_2(2), operand_2(2) => 
                           operand_2(1), operand_2(1) => operand_2(0), p(32) =>
                           p_31_port, p(31) => p_30_port, p(30) => p_29_port, 
                           p(29) => p_28_port, p(28) => p_27_port, p(27) => 
                           p_26_port, p(26) => p_25_port, p(25) => p_24_port, 
                           p(24) => p_23_port, p(23) => p_22_port, p(22) => 
                           p_21_port, p(21) => p_20_port, p(20) => p_19_port, 
                           p(19) => p_18_port, p(18) => p_17_port, p(17) => 
                           p_16_port, p(16) => p_15_port, p(15) => p_14_port, 
                           p(14) => p_13_port, p(13) => p_12_port, p(12) => 
                           p_11_port, p(11) => p_10_port, p(10) => p_9_port, 
                           p(9) => p_8_port, p(8) => p_7_port, p(7) => p_6_port
                           , p(6) => p_5_port, p(5) => p_4_port, p(4) => 
                           p_3_port, p(3) => p_2_port, p(2) => p_1_port, p(1) 
                           => p_0_port, g(32) => g_31_port, g(31) => g_30_port,
                           g(30) => g_29_port, g(29) => g_28_port, g(28) => 
                           g_27_port, g(27) => g_26_port, g(26) => g_25_port, 
                           g(25) => g_24_port, g(24) => g_23_port, g(23) => 
                           g_22_port, g(22) => g_21_port, g(21) => g_20_port, 
                           g(20) => g_19_port, g(19) => g_18_port, g(18) => 
                           g_17_port, g(17) => g_16_port, g(16) => g_15_port, 
                           g(15) => g_14_port, g(14) => g_13_port, g(13) => 
                           g_12_port, g(12) => g_11_port, g(11) => g_10_port, 
                           g(10) => g_9_port, g(9) => g_8_port, g(8) => 
                           g_7_port, g(7) => g_6_port, g(6) => g_5_port, g(5) 
                           => g_4_port, g(4) => g_3_port, g(3) => g_2_port, 
                           g(2) => g_1_port, g(1) => g_0_port);
   flgblock : g_block_carry port map( Gik => g_1_port, Pik => p_1_port, Gk1j =>
                           g_0_port, Pk1j => p_0_port, carry_in => carry_in, 
                           Gij => g_matrix_0_0_port);
   flpgblock_1 : pg_block_0 port map( Gik => g_3_port, Pik => p_3_port, Gk1j =>
                           g_2_port, Pk1j => p_2_port, Gij => g_matrix_0_1_port
                           , Pij => p_matrix_0_1_port);
   flpgblock_2 : pg_block_26 port map( Gik => g_5_port, Pik => p_5_port, Gk1j 
                           => g_4_port, Pk1j => p_4_port, Gij => 
                           g_matrix_0_2_port, Pij => p_matrix_0_2_port);
   flpgblock_3 : pg_block_25 port map( Gik => g_7_port, Pik => p_7_port, Gk1j 
                           => g_6_port, Pk1j => p_6_port, Gij => 
                           g_matrix_0_3_port, Pij => p_matrix_0_3_port);
   flpgblock_4 : pg_block_24 port map( Gik => g_9_port, Pik => p_9_port, Gk1j 
                           => g_8_port, Pk1j => p_8_port, Gij => 
                           g_matrix_0_4_port, Pij => p_matrix_0_4_port);
   flpgblock_5 : pg_block_23 port map( Gik => g_11_port, Pik => p_11_port, Gk1j
                           => g_10_port, Pk1j => p_10_port, Gij => 
                           g_matrix_0_5_port, Pij => p_matrix_0_5_port);
   flpgblock_6 : pg_block_22 port map( Gik => g_13_port, Pik => p_13_port, Gk1j
                           => g_12_port, Pk1j => p_12_port, Gij => 
                           g_matrix_0_6_port, Pij => p_matrix_0_6_port);
   flpgblock_7 : pg_block_21 port map( Gik => g_15_port, Pik => p_15_port, Gk1j
                           => g_14_port, Pk1j => p_14_port, Gij => 
                           g_matrix_0_7_port, Pij => p_matrix_0_7_port);
   flpgblock_8 : pg_block_20 port map( Gik => g_17_port, Pik => p_17_port, Gk1j
                           => g_16_port, Pk1j => p_16_port, Gij => 
                           g_matrix_0_8_port, Pij => p_matrix_0_8_port);
   flpgblock_9 : pg_block_19 port map( Gik => g_19_port, Pik => p_19_port, Gk1j
                           => g_18_port, Pk1j => p_18_port, Gij => 
                           g_matrix_0_9_port, Pij => p_matrix_0_9_port);
   flpgblock_10 : pg_block_18 port map( Gik => g_21_port, Pik => p_21_port, 
                           Gk1j => g_20_port, Pk1j => p_20_port, Gij => 
                           g_matrix_0_10_port, Pij => p_matrix_0_10_port);
   flpgblock_11 : pg_block_17 port map( Gik => g_23_port, Pik => p_23_port, 
                           Gk1j => g_22_port, Pk1j => p_22_port, Gij => 
                           g_matrix_0_11_port, Pij => p_matrix_0_11_port);
   flpgblock_12 : pg_block_16 port map( Gik => g_25_port, Pik => p_25_port, 
                           Gk1j => g_24_port, Pk1j => p_24_port, Gij => 
                           g_matrix_0_12_port, Pij => p_matrix_0_12_port);
   flpgblock_13 : pg_block_15 port map( Gik => g_27_port, Pik => p_27_port, 
                           Gk1j => g_26_port, Pk1j => p_26_port, Gij => 
                           g_matrix_0_13_port, Pij => p_matrix_0_13_port);
   flpgblock_14 : pg_block_14 port map( Gik => g_29_port, Pik => p_29_port, 
                           Gk1j => g_28_port, Pk1j => p_28_port, Gij => 
                           g_matrix_0_14_port, Pij => p_matrix_0_14_port);
   flpgblock_15 : pg_block_13 port map( Gik => g_31_port, Pik => p_31_port, 
                           Gk1j => g_30_port, Pk1j => p_30_port, Gij => 
                           g_matrix_0_15_port, Pij => p_matrix_0_15_port);
   slgblock : g_block_0 port map( Gik => g_matrix_0_1_port, Pik => 
                           p_matrix_0_1_port, Gk1j => g_matrix_0_0_port, Gij =>
                           carry_out_0_port);
   slpgblock_1 : pg_block_12 port map( Gik => g_matrix_0_3_port, Pik => 
                           p_matrix_0_3_port, Gk1j => g_matrix_0_2_port, Pk1j 
                           => p_matrix_0_2_port, Gij => g_matrix_1_1_port, Pij 
                           => p_matrix_1_1_port);
   slpgblock_2 : pg_block_11 port map( Gik => g_matrix_0_5_port, Pik => 
                           p_matrix_0_5_port, Gk1j => g_matrix_0_4_port, Pk1j 
                           => p_matrix_0_4_port, Gij => g_matrix_1_2_port, Pij 
                           => p_matrix_1_2_port);
   slpgblock_3 : pg_block_10 port map( Gik => g_matrix_0_7_port, Pik => 
                           p_matrix_0_7_port, Gk1j => g_matrix_0_6_port, Pk1j 
                           => p_matrix_0_6_port, Gij => g_matrix_1_3_port, Pij 
                           => p_matrix_1_3_port);
   slpgblock_4 : pg_block_9 port map( Gik => g_matrix_0_9_port, Pik => 
                           p_matrix_0_9_port, Gk1j => g_matrix_0_8_port, Pk1j 
                           => p_matrix_0_8_port, Gij => g_matrix_1_4_port, Pij 
                           => p_matrix_1_4_port);
   slpgblock_5 : pg_block_8 port map( Gik => g_matrix_0_11_port, Pik => 
                           p_matrix_0_11_port, Gk1j => g_matrix_0_10_port, Pk1j
                           => p_matrix_0_10_port, Gij => g_matrix_1_5_port, Pij
                           => p_matrix_1_5_port);
   slpgblock_6 : pg_block_7 port map( Gik => g_matrix_0_13_port, Pik => 
                           p_matrix_0_13_port, Gk1j => g_matrix_0_12_port, Pk1j
                           => p_matrix_0_12_port, Gij => g_matrix_1_6_port, Pij
                           => p_matrix_1_6_port);
   slpgblock_7 : pg_block_6 port map( Gik => g_matrix_0_15_port, Pik => 
                           p_matrix_0_15_port, Gk1j => g_matrix_0_14_port, Pk1j
                           => p_matrix_0_14_port, Gij => g_matrix_1_7_port, Pij
                           => p_matrix_1_7_port);
   olgblock_2_1 : g_block_7 port map( Gik => g_matrix_1_1_port, Pik => 
                           p_matrix_1_1_port, Gk1j => carry_out_0_port, Gij => 
                           carry_out_1_port);
   olpgblock_2_3 : pg_block_5 port map( Gik => g_matrix_1_3_port, Pik => 
                           p_matrix_1_3_port, Gk1j => g_matrix_1_1_port, Pk1j 
                           => p_matrix_1_1_port, Gij => g_matrix_2_3_port, Pij 
                           => p_matrix_2_3_port);
   olpgblock_2_5 : pg_block_4 port map( Gik => g_matrix_1_5_port, Pik => 
                           p_matrix_1_5_port, Gk1j => g_matrix_1_3_port, Pk1j 
                           => p_matrix_1_3_port, Gij => g_matrix_2_5_port, Pij 
                           => p_matrix_2_5_port);
   olpgblock_2_7 : pg_block_3 port map( Gik => g_matrix_1_7_port, Pik => 
                           p_matrix_1_7_port, Gk1j => g_matrix_1_5_port, Pk1j 
                           => p_matrix_1_5_port, Gij => g_matrix_2_7_port, Pij 
                           => p_matrix_2_7_port);
   olgblock_3_2 : g_block_6 port map( Gik => g_matrix_1_2_port, Pik => 
                           p_matrix_1_2_port, Gk1j => carry_out_1_port, Gij => 
                           carry_out_2_port);
   olgblock_3_3 : g_block_5 port map( Gik => g_matrix_2_3_port, Pik => 
                           p_matrix_2_3_port, Gk1j => carry_out_1_port, Gij => 
                           carry_out_3_port);
   olpgblock_3_6 : pg_block_2 port map( Gik => g_matrix_1_6_port, Pik => 
                           p_matrix_1_6_port, Gk1j => g_matrix_1_4_port, Pk1j 
                           => p_matrix_1_4_port, Gij => g_matrix_3_6_port, Pij 
                           => p_matrix_3_6_port);
   olpgblock_3_7 : pg_block_1 port map( Gik => g_matrix_2_7_port, Pik => 
                           p_matrix_2_7_port, Gk1j => g_matrix_2_5_port, Pk1j 
                           => p_matrix_2_5_port, Gij => g_matrix_3_7_port, Pij 
                           => p_matrix_3_7_port);
   olgblock_4_4 : g_block_4 port map( Gik => g_matrix_1_4_port, Pik => 
                           p_matrix_1_4_port, Gk1j => carry_out_2_port, Gij => 
                           carry_out_4_port);
   olgblock_4_5 : g_block_3 port map( Gik => g_matrix_2_5_port, Pik => 
                           p_matrix_2_5_port, Gk1j => carry_out_2_port, Gij => 
                           carry_out_5_port);
   olgblock_4_6 : g_block_2 port map( Gik => g_matrix_3_6_port, Pik => 
                           p_matrix_3_6_port, Gk1j => carry_out_2_port, Gij => 
                           carry_out_6_port);
   olgblock_4_7 : g_block_1 port map( Gik => g_matrix_3_7_port, Pik => 
                           p_matrix_3_7_port, Gk1j => carry_out_2_port, Gij => 
                           carry_out_7_port);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shifter_nbit32 is

   port( r1, r2 : in std_logic_vector (31 downto 0);  conf : in 
         std_logic_vector (1 downto 0);  shifted_out : out std_logic_vector (31
         downto 0));

end shifter_nbit32;

architecture SYN_structural of shifter_nbit32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX81_N32
      port( a, b, c, d, e, f, g, h : in std_logic_vector (31 downto 0);  sel : 
            in std_logic_vector (2 downto 0);  y : out std_logic_vector (31 
            downto 0));
   end component;
   
   component MUX41_N40
      port( a, b, c, d : in std_logic_vector (39 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  y : out std_logic_vector (39 downto
            0));
   end component;
   
   component MUX21_N40_1
      port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (39 downto 0));
   end component;
   
   component MUX21_N40_2
      port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (39 downto 0));
   end component;
   
   component MUX21_N40_3
      port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (39 downto 0));
   end component;
   
   component MUX21_N40_0
      port( a, b : in std_logic_vector (39 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (39 downto 0));
   end component;
   
   signal X_Logic0_port, right_first_level_3_39_port, 
      final_first_level_0_39_port, final_first_level_0_38_port, 
      final_first_level_0_37_port, final_first_level_0_36_port, 
      final_first_level_0_35_port, final_first_level_0_34_port, 
      final_first_level_0_33_port, final_first_level_0_32_port, 
      final_first_level_0_31_port, final_first_level_0_30_port, 
      final_first_level_0_29_port, final_first_level_0_28_port, 
      final_first_level_0_27_port, final_first_level_0_26_port, 
      final_first_level_0_25_port, final_first_level_0_24_port, 
      final_first_level_0_23_port, final_first_level_0_22_port, 
      final_first_level_0_21_port, final_first_level_0_20_port, 
      final_first_level_0_19_port, final_first_level_0_18_port, 
      final_first_level_0_17_port, final_first_level_0_16_port, 
      final_first_level_0_15_port, final_first_level_0_14_port, 
      final_first_level_0_13_port, final_first_level_0_12_port, 
      final_first_level_0_11_port, final_first_level_0_10_port, 
      final_first_level_0_9_port, final_first_level_0_8_port, 
      final_first_level_0_7_port, final_first_level_0_6_port, 
      final_first_level_0_5_port, final_first_level_0_4_port, 
      final_first_level_0_3_port, final_first_level_0_2_port, 
      final_first_level_0_1_port, final_first_level_0_0_port, 
      final_first_level_1_39_port, final_first_level_1_38_port, 
      final_first_level_1_37_port, final_first_level_1_36_port, 
      final_first_level_1_35_port, final_first_level_1_34_port, 
      final_first_level_1_33_port, final_first_level_1_32_port, 
      final_first_level_1_31_port, final_first_level_1_30_port, 
      final_first_level_1_29_port, final_first_level_1_28_port, 
      final_first_level_1_27_port, final_first_level_1_26_port, 
      final_first_level_1_25_port, final_first_level_1_24_port, 
      final_first_level_1_23_port, final_first_level_1_22_port, 
      final_first_level_1_21_port, final_first_level_1_20_port, 
      final_first_level_1_19_port, final_first_level_1_18_port, 
      final_first_level_1_17_port, final_first_level_1_16_port, 
      final_first_level_1_15_port, final_first_level_1_14_port, 
      final_first_level_1_13_port, final_first_level_1_12_port, 
      final_first_level_1_11_port, final_first_level_1_10_port, 
      final_first_level_1_9_port, final_first_level_1_8_port, 
      final_first_level_1_7_port, final_first_level_1_6_port, 
      final_first_level_1_5_port, final_first_level_1_4_port, 
      final_first_level_1_3_port, final_first_level_1_2_port, 
      final_first_level_1_1_port, final_first_level_1_0_port, 
      final_first_level_2_39_port, final_first_level_2_38_port, 
      final_first_level_2_37_port, final_first_level_2_36_port, 
      final_first_level_2_35_port, final_first_level_2_34_port, 
      final_first_level_2_33_port, final_first_level_2_32_port, 
      final_first_level_2_31_port, final_first_level_2_30_port, 
      final_first_level_2_29_port, final_first_level_2_28_port, 
      final_first_level_2_27_port, final_first_level_2_26_port, 
      final_first_level_2_25_port, final_first_level_2_24_port, 
      final_first_level_2_23_port, final_first_level_2_22_port, 
      final_first_level_2_21_port, final_first_level_2_20_port, 
      final_first_level_2_19_port, final_first_level_2_18_port, 
      final_first_level_2_17_port, final_first_level_2_16_port, 
      final_first_level_2_15_port, final_first_level_2_14_port, 
      final_first_level_2_13_port, final_first_level_2_12_port, 
      final_first_level_2_11_port, final_first_level_2_10_port, 
      final_first_level_2_9_port, final_first_level_2_8_port, 
      final_first_level_2_7_port, final_first_level_2_6_port, 
      final_first_level_2_5_port, final_first_level_2_4_port, 
      final_first_level_2_3_port, final_first_level_2_2_port, 
      final_first_level_2_1_port, final_first_level_2_0_port, 
      final_first_level_3_39_port, final_first_level_3_38_port, 
      final_first_level_3_37_port, final_first_level_3_36_port, 
      final_first_level_3_35_port, final_first_level_3_34_port, 
      final_first_level_3_33_port, final_first_level_3_32_port, 
      final_first_level_3_31_port, final_first_level_3_30_port, 
      final_first_level_3_29_port, final_first_level_3_28_port, 
      final_first_level_3_27_port, final_first_level_3_26_port, 
      final_first_level_3_25_port, final_first_level_3_24_port, 
      final_first_level_3_23_port, final_first_level_3_22_port, 
      final_first_level_3_21_port, final_first_level_3_20_port, 
      final_first_level_3_19_port, final_first_level_3_18_port, 
      final_first_level_3_17_port, final_first_level_3_16_port, 
      final_first_level_3_15_port, final_first_level_3_14_port, 
      final_first_level_3_13_port, final_first_level_3_12_port, 
      final_first_level_3_11_port, final_first_level_3_10_port, 
      final_first_level_3_9_port, final_first_level_3_8_port, 
      final_first_level_3_7_port, final_first_level_3_6_port, 
      final_first_level_3_5_port, final_first_level_3_4_port, 
      final_first_level_3_3_port, final_first_level_3_2_port, 
      final_first_level_3_1_port, final_first_level_3_0_port, 
      final_first_level_mask_38_port, final_first_level_mask_37_port, 
      final_first_level_mask_36_port, final_first_level_mask_35_port, 
      final_first_level_mask_34_port, final_first_level_mask_33_port, 
      final_first_level_mask_32_port, final_first_level_mask_31_port, 
      final_first_level_mask_30_port, final_first_level_mask_29_port, 
      final_first_level_mask_28_port, final_first_level_mask_27_port, 
      final_first_level_mask_26_port, final_first_level_mask_25_port, 
      final_first_level_mask_24_port, final_first_level_mask_23_port, 
      final_first_level_mask_22_port, final_first_level_mask_21_port, 
      final_first_level_mask_20_port, final_first_level_mask_19_port, 
      final_first_level_mask_18_port, final_first_level_mask_17_port, 
      final_first_level_mask_16_port, final_first_level_mask_15_port, 
      final_first_level_mask_14_port, final_first_level_mask_13_port, 
      final_first_level_mask_12_port, final_first_level_mask_11_port, 
      final_first_level_mask_10_port, final_first_level_mask_9_port, 
      final_first_level_mask_8_port, final_first_level_mask_7_port, 
      final_first_level_mask_6_port, final_first_level_mask_5_port, 
      final_first_level_mask_4_port, final_first_level_mask_3_port, 
      final_first_level_mask_2_port, final_first_level_mask_1_port, 
      final_first_level_mask_0_port, third_level_sel_2_port, 
      third_level_sel_1_port, third_level_sel_0_port, n_1163 : std_logic;

begin
   
   X_Logic0_port <= '0';
   MUX21_i_1 : MUX21_N40_0 port map( a(39) => right_first_level_3_39_port, 
                           a(38) => right_first_level_3_39_port, a(37) => 
                           right_first_level_3_39_port, a(36) => 
                           right_first_level_3_39_port, a(35) => 
                           right_first_level_3_39_port, a(34) => 
                           right_first_level_3_39_port, a(33) => 
                           right_first_level_3_39_port, a(32) => 
                           right_first_level_3_39_port, a(31) => r1(31), a(30) 
                           => r1(30), a(29) => r1(29), a(28) => r1(28), a(27) 
                           => r1(27), a(26) => r1(26), a(25) => r1(25), a(24) 
                           => r1(24), a(23) => r1(23), a(22) => r1(22), a(21) 
                           => r1(21), a(20) => r1(20), a(19) => r1(19), a(18) 
                           => r1(18), a(17) => r1(17), a(16) => r1(16), a(15) 
                           => r1(15), a(14) => r1(14), a(13) => r1(13), a(12) 
                           => r1(12), a(11) => r1(11), a(10) => r1(10), a(9) =>
                           r1(9), a(8) => r1(8), a(7) => r1(7), a(6) => r1(6), 
                           a(5) => r1(5), a(4) => r1(4), a(3) => r1(3), a(2) =>
                           r1(2), a(1) => r1(1), a(0) => r1(0), b(39) => 
                           X_Logic0_port, b(38) => r1(31), b(37) => r1(30), 
                           b(36) => r1(29), b(35) => r1(28), b(34) => r1(27), 
                           b(33) => r1(26), b(32) => r1(25), b(31) => r1(24), 
                           b(30) => r1(23), b(29) => r1(22), b(28) => r1(21), 
                           b(27) => r1(20), b(26) => r1(19), b(25) => r1(18), 
                           b(24) => r1(17), b(23) => r1(16), b(22) => r1(15), 
                           b(21) => r1(14), b(20) => r1(13), b(19) => r1(12), 
                           b(18) => r1(11), b(17) => r1(10), b(16) => r1(9), 
                           b(15) => r1(8), b(14) => r1(7), b(13) => r1(6), 
                           b(12) => r1(5), b(11) => r1(4), b(10) => r1(3), b(9)
                           => r1(2), b(8) => r1(1), b(7) => r1(0), b(6) => 
                           X_Logic0_port, b(5) => X_Logic0_port, b(4) => 
                           X_Logic0_port, b(3) => X_Logic0_port, b(2) => 
                           X_Logic0_port, b(1) => X_Logic0_port, b(0) => 
                           X_Logic0_port, sel => conf(0), y(39) => 
                           final_first_level_0_39_port, y(38) => 
                           final_first_level_0_38_port, y(37) => 
                           final_first_level_0_37_port, y(36) => 
                           final_first_level_0_36_port, y(35) => 
                           final_first_level_0_35_port, y(34) => 
                           final_first_level_0_34_port, y(33) => 
                           final_first_level_0_33_port, y(32) => 
                           final_first_level_0_32_port, y(31) => 
                           final_first_level_0_31_port, y(30) => 
                           final_first_level_0_30_port, y(29) => 
                           final_first_level_0_29_port, y(28) => 
                           final_first_level_0_28_port, y(27) => 
                           final_first_level_0_27_port, y(26) => 
                           final_first_level_0_26_port, y(25) => 
                           final_first_level_0_25_port, y(24) => 
                           final_first_level_0_24_port, y(23) => 
                           final_first_level_0_23_port, y(22) => 
                           final_first_level_0_22_port, y(21) => 
                           final_first_level_0_21_port, y(20) => 
                           final_first_level_0_20_port, y(19) => 
                           final_first_level_0_19_port, y(18) => 
                           final_first_level_0_18_port, y(17) => 
                           final_first_level_0_17_port, y(16) => 
                           final_first_level_0_16_port, y(15) => 
                           final_first_level_0_15_port, y(14) => 
                           final_first_level_0_14_port, y(13) => 
                           final_first_level_0_13_port, y(12) => 
                           final_first_level_0_12_port, y(11) => 
                           final_first_level_0_11_port, y(10) => 
                           final_first_level_0_10_port, y(9) => 
                           final_first_level_0_9_port, y(8) => 
                           final_first_level_0_8_port, y(7) => 
                           final_first_level_0_7_port, y(6) => 
                           final_first_level_0_6_port, y(5) => 
                           final_first_level_0_5_port, y(4) => 
                           final_first_level_0_4_port, y(3) => 
                           final_first_level_0_3_port, y(2) => 
                           final_first_level_0_2_port, y(1) => 
                           final_first_level_0_1_port, y(0) => 
                           final_first_level_0_0_port);
   MUX21_i_2 : MUX21_N40_3 port map( a(39) => right_first_level_3_39_port, 
                           a(38) => right_first_level_3_39_port, a(37) => 
                           right_first_level_3_39_port, a(36) => 
                           right_first_level_3_39_port, a(35) => 
                           right_first_level_3_39_port, a(34) => 
                           right_first_level_3_39_port, a(33) => 
                           right_first_level_3_39_port, a(32) => 
                           right_first_level_3_39_port, a(31) => 
                           right_first_level_3_39_port, a(30) => 
                           right_first_level_3_39_port, a(29) => 
                           right_first_level_3_39_port, a(28) => 
                           right_first_level_3_39_port, a(27) => 
                           right_first_level_3_39_port, a(26) => 
                           right_first_level_3_39_port, a(25) => 
                           right_first_level_3_39_port, a(24) => 
                           right_first_level_3_39_port, a(23) => r1(31), a(22) 
                           => r1(30), a(21) => r1(29), a(20) => r1(28), a(19) 
                           => r1(27), a(18) => r1(26), a(17) => r1(25), a(16) 
                           => r1(24), a(15) => r1(23), a(14) => r1(22), a(13) 
                           => r1(21), a(12) => r1(20), a(11) => r1(19), a(10) 
                           => r1(18), a(9) => r1(17), a(8) => r1(16), a(7) => 
                           r1(15), a(6) => r1(14), a(5) => r1(13), a(4) => 
                           r1(12), a(3) => r1(11), a(2) => r1(10), a(1) => 
                           r1(9), a(0) => r1(8), b(39) => X_Logic0_port, b(38) 
                           => r1(23), b(37) => r1(22), b(36) => r1(21), b(35) 
                           => r1(20), b(34) => r1(19), b(33) => r1(18), b(32) 
                           => r1(17), b(31) => r1(16), b(30) => r1(15), b(29) 
                           => r1(14), b(28) => r1(13), b(27) => r1(12), b(26) 
                           => r1(11), b(25) => r1(10), b(24) => r1(9), b(23) =>
                           r1(8), b(22) => r1(7), b(21) => r1(6), b(20) => 
                           r1(5), b(19) => r1(4), b(18) => r1(3), b(17) => 
                           r1(2), b(16) => r1(1), b(15) => r1(0), b(14) => 
                           X_Logic0_port, b(13) => X_Logic0_port, b(12) => 
                           X_Logic0_port, b(11) => X_Logic0_port, b(10) => 
                           X_Logic0_port, b(9) => X_Logic0_port, b(8) => 
                           X_Logic0_port, b(7) => X_Logic0_port, b(6) => 
                           X_Logic0_port, b(5) => X_Logic0_port, b(4) => 
                           X_Logic0_port, b(3) => X_Logic0_port, b(2) => 
                           X_Logic0_port, b(1) => X_Logic0_port, b(0) => 
                           X_Logic0_port, sel => conf(0), y(39) => 
                           final_first_level_1_39_port, y(38) => 
                           final_first_level_1_38_port, y(37) => 
                           final_first_level_1_37_port, y(36) => 
                           final_first_level_1_36_port, y(35) => 
                           final_first_level_1_35_port, y(34) => 
                           final_first_level_1_34_port, y(33) => 
                           final_first_level_1_33_port, y(32) => 
                           final_first_level_1_32_port, y(31) => 
                           final_first_level_1_31_port, y(30) => 
                           final_first_level_1_30_port, y(29) => 
                           final_first_level_1_29_port, y(28) => 
                           final_first_level_1_28_port, y(27) => 
                           final_first_level_1_27_port, y(26) => 
                           final_first_level_1_26_port, y(25) => 
                           final_first_level_1_25_port, y(24) => 
                           final_first_level_1_24_port, y(23) => 
                           final_first_level_1_23_port, y(22) => 
                           final_first_level_1_22_port, y(21) => 
                           final_first_level_1_21_port, y(20) => 
                           final_first_level_1_20_port, y(19) => 
                           final_first_level_1_19_port, y(18) => 
                           final_first_level_1_18_port, y(17) => 
                           final_first_level_1_17_port, y(16) => 
                           final_first_level_1_16_port, y(15) => 
                           final_first_level_1_15_port, y(14) => 
                           final_first_level_1_14_port, y(13) => 
                           final_first_level_1_13_port, y(12) => 
                           final_first_level_1_12_port, y(11) => 
                           final_first_level_1_11_port, y(10) => 
                           final_first_level_1_10_port, y(9) => 
                           final_first_level_1_9_port, y(8) => 
                           final_first_level_1_8_port, y(7) => 
                           final_first_level_1_7_port, y(6) => 
                           final_first_level_1_6_port, y(5) => 
                           final_first_level_1_5_port, y(4) => 
                           final_first_level_1_4_port, y(3) => 
                           final_first_level_1_3_port, y(2) => 
                           final_first_level_1_2_port, y(1) => 
                           final_first_level_1_1_port, y(0) => 
                           final_first_level_1_0_port);
   MUX21_i_3 : MUX21_N40_2 port map( a(39) => right_first_level_3_39_port, 
                           a(38) => right_first_level_3_39_port, a(37) => 
                           right_first_level_3_39_port, a(36) => 
                           right_first_level_3_39_port, a(35) => 
                           right_first_level_3_39_port, a(34) => 
                           right_first_level_3_39_port, a(33) => 
                           right_first_level_3_39_port, a(32) => 
                           right_first_level_3_39_port, a(31) => 
                           right_first_level_3_39_port, a(30) => 
                           right_first_level_3_39_port, a(29) => 
                           right_first_level_3_39_port, a(28) => 
                           right_first_level_3_39_port, a(27) => 
                           right_first_level_3_39_port, a(26) => 
                           right_first_level_3_39_port, a(25) => 
                           right_first_level_3_39_port, a(24) => 
                           right_first_level_3_39_port, a(23) => 
                           right_first_level_3_39_port, a(22) => 
                           right_first_level_3_39_port, a(21) => 
                           right_first_level_3_39_port, a(20) => 
                           right_first_level_3_39_port, a(19) => 
                           right_first_level_3_39_port, a(18) => 
                           right_first_level_3_39_port, a(17) => 
                           right_first_level_3_39_port, a(16) => 
                           right_first_level_3_39_port, a(15) => r1(31), a(14) 
                           => r1(30), a(13) => r1(29), a(12) => r1(28), a(11) 
                           => r1(27), a(10) => r1(26), a(9) => r1(25), a(8) => 
                           r1(24), a(7) => r1(23), a(6) => r1(22), a(5) => 
                           r1(21), a(4) => r1(20), a(3) => r1(19), a(2) => 
                           r1(18), a(1) => r1(17), a(0) => r1(16), b(39) => 
                           X_Logic0_port, b(38) => r1(15), b(37) => r1(14), 
                           b(36) => r1(13), b(35) => r1(12), b(34) => r1(11), 
                           b(33) => r1(10), b(32) => r1(9), b(31) => r1(8), 
                           b(30) => r1(7), b(29) => r1(6), b(28) => r1(5), 
                           b(27) => r1(4), b(26) => r1(3), b(25) => r1(2), 
                           b(24) => r1(1), b(23) => r1(0), b(22) => 
                           X_Logic0_port, b(21) => X_Logic0_port, b(20) => 
                           X_Logic0_port, b(19) => X_Logic0_port, b(18) => 
                           X_Logic0_port, b(17) => X_Logic0_port, b(16) => 
                           X_Logic0_port, b(15) => X_Logic0_port, b(14) => 
                           X_Logic0_port, b(13) => X_Logic0_port, b(12) => 
                           X_Logic0_port, b(11) => X_Logic0_port, b(10) => 
                           X_Logic0_port, b(9) => X_Logic0_port, b(8) => 
                           X_Logic0_port, b(7) => X_Logic0_port, b(6) => 
                           X_Logic0_port, b(5) => X_Logic0_port, b(4) => 
                           X_Logic0_port, b(3) => X_Logic0_port, b(2) => 
                           X_Logic0_port, b(1) => X_Logic0_port, b(0) => 
                           X_Logic0_port, sel => conf(0), y(39) => 
                           final_first_level_2_39_port, y(38) => 
                           final_first_level_2_38_port, y(37) => 
                           final_first_level_2_37_port, y(36) => 
                           final_first_level_2_36_port, y(35) => 
                           final_first_level_2_35_port, y(34) => 
                           final_first_level_2_34_port, y(33) => 
                           final_first_level_2_33_port, y(32) => 
                           final_first_level_2_32_port, y(31) => 
                           final_first_level_2_31_port, y(30) => 
                           final_first_level_2_30_port, y(29) => 
                           final_first_level_2_29_port, y(28) => 
                           final_first_level_2_28_port, y(27) => 
                           final_first_level_2_27_port, y(26) => 
                           final_first_level_2_26_port, y(25) => 
                           final_first_level_2_25_port, y(24) => 
                           final_first_level_2_24_port, y(23) => 
                           final_first_level_2_23_port, y(22) => 
                           final_first_level_2_22_port, y(21) => 
                           final_first_level_2_21_port, y(20) => 
                           final_first_level_2_20_port, y(19) => 
                           final_first_level_2_19_port, y(18) => 
                           final_first_level_2_18_port, y(17) => 
                           final_first_level_2_17_port, y(16) => 
                           final_first_level_2_16_port, y(15) => 
                           final_first_level_2_15_port, y(14) => 
                           final_first_level_2_14_port, y(13) => 
                           final_first_level_2_13_port, y(12) => 
                           final_first_level_2_12_port, y(11) => 
                           final_first_level_2_11_port, y(10) => 
                           final_first_level_2_10_port, y(9) => 
                           final_first_level_2_9_port, y(8) => 
                           final_first_level_2_8_port, y(7) => 
                           final_first_level_2_7_port, y(6) => 
                           final_first_level_2_6_port, y(5) => 
                           final_first_level_2_5_port, y(4) => 
                           final_first_level_2_4_port, y(3) => 
                           final_first_level_2_3_port, y(2) => 
                           final_first_level_2_2_port, y(1) => 
                           final_first_level_2_1_port, y(0) => 
                           final_first_level_2_0_port);
   MUX21_i_4 : MUX21_N40_1 port map( a(39) => right_first_level_3_39_port, 
                           a(38) => right_first_level_3_39_port, a(37) => 
                           right_first_level_3_39_port, a(36) => 
                           right_first_level_3_39_port, a(35) => 
                           right_first_level_3_39_port, a(34) => 
                           right_first_level_3_39_port, a(33) => 
                           right_first_level_3_39_port, a(32) => 
                           right_first_level_3_39_port, a(31) => 
                           right_first_level_3_39_port, a(30) => 
                           right_first_level_3_39_port, a(29) => 
                           right_first_level_3_39_port, a(28) => 
                           right_first_level_3_39_port, a(27) => 
                           right_first_level_3_39_port, a(26) => 
                           right_first_level_3_39_port, a(25) => 
                           right_first_level_3_39_port, a(24) => 
                           right_first_level_3_39_port, a(23) => 
                           right_first_level_3_39_port, a(22) => 
                           right_first_level_3_39_port, a(21) => 
                           right_first_level_3_39_port, a(20) => 
                           right_first_level_3_39_port, a(19) => 
                           right_first_level_3_39_port, a(18) => 
                           right_first_level_3_39_port, a(17) => 
                           right_first_level_3_39_port, a(16) => 
                           right_first_level_3_39_port, a(15) => 
                           right_first_level_3_39_port, a(14) => 
                           right_first_level_3_39_port, a(13) => 
                           right_first_level_3_39_port, a(12) => 
                           right_first_level_3_39_port, a(11) => 
                           right_first_level_3_39_port, a(10) => 
                           right_first_level_3_39_port, a(9) => 
                           right_first_level_3_39_port, a(8) => 
                           right_first_level_3_39_port, a(7) => r1(31), a(6) =>
                           r1(30), a(5) => r1(29), a(4) => r1(28), a(3) => 
                           r1(27), a(2) => r1(26), a(1) => r1(25), a(0) => 
                           r1(24), b(39) => X_Logic0_port, b(38) => r1(7), 
                           b(37) => r1(6), b(36) => r1(5), b(35) => r1(4), 
                           b(34) => r1(3), b(33) => r1(2), b(32) => r1(1), 
                           b(31) => r1(0), b(30) => X_Logic0_port, b(29) => 
                           X_Logic0_port, b(28) => X_Logic0_port, b(27) => 
                           X_Logic0_port, b(26) => X_Logic0_port, b(25) => 
                           X_Logic0_port, b(24) => X_Logic0_port, b(23) => 
                           X_Logic0_port, b(22) => X_Logic0_port, b(21) => 
                           X_Logic0_port, b(20) => X_Logic0_port, b(19) => 
                           X_Logic0_port, b(18) => X_Logic0_port, b(17) => 
                           X_Logic0_port, b(16) => X_Logic0_port, b(15) => 
                           X_Logic0_port, b(14) => X_Logic0_port, b(13) => 
                           X_Logic0_port, b(12) => X_Logic0_port, b(11) => 
                           X_Logic0_port, b(10) => X_Logic0_port, b(9) => 
                           X_Logic0_port, b(8) => X_Logic0_port, b(7) => 
                           X_Logic0_port, b(6) => X_Logic0_port, b(5) => 
                           X_Logic0_port, b(4) => X_Logic0_port, b(3) => 
                           X_Logic0_port, b(2) => X_Logic0_port, b(1) => 
                           X_Logic0_port, b(0) => X_Logic0_port, sel => conf(0)
                           , y(39) => final_first_level_3_39_port, y(38) => 
                           final_first_level_3_38_port, y(37) => 
                           final_first_level_3_37_port, y(36) => 
                           final_first_level_3_36_port, y(35) => 
                           final_first_level_3_35_port, y(34) => 
                           final_first_level_3_34_port, y(33) => 
                           final_first_level_3_33_port, y(32) => 
                           final_first_level_3_32_port, y(31) => 
                           final_first_level_3_31_port, y(30) => 
                           final_first_level_3_30_port, y(29) => 
                           final_first_level_3_29_port, y(28) => 
                           final_first_level_3_28_port, y(27) => 
                           final_first_level_3_27_port, y(26) => 
                           final_first_level_3_26_port, y(25) => 
                           final_first_level_3_25_port, y(24) => 
                           final_first_level_3_24_port, y(23) => 
                           final_first_level_3_23_port, y(22) => 
                           final_first_level_3_22_port, y(21) => 
                           final_first_level_3_21_port, y(20) => 
                           final_first_level_3_20_port, y(19) => 
                           final_first_level_3_19_port, y(18) => 
                           final_first_level_3_18_port, y(17) => 
                           final_first_level_3_17_port, y(16) => 
                           final_first_level_3_16_port, y(15) => 
                           final_first_level_3_15_port, y(14) => 
                           final_first_level_3_14_port, y(13) => 
                           final_first_level_3_13_port, y(12) => 
                           final_first_level_3_12_port, y(11) => 
                           final_first_level_3_11_port, y(10) => 
                           final_first_level_3_10_port, y(9) => 
                           final_first_level_3_9_port, y(8) => 
                           final_first_level_3_8_port, y(7) => 
                           final_first_level_3_7_port, y(6) => 
                           final_first_level_3_6_port, y(5) => 
                           final_first_level_3_5_port, y(4) => 
                           final_first_level_3_4_port, y(3) => 
                           final_first_level_3_3_port, y(2) => 
                           final_first_level_3_2_port, y(1) => 
                           final_first_level_3_1_port, y(0) => 
                           final_first_level_3_0_port);
   MUX41_level_2 : MUX41_N40 port map( a(39) => final_first_level_0_39_port, 
                           a(38) => final_first_level_0_38_port, a(37) => 
                           final_first_level_0_37_port, a(36) => 
                           final_first_level_0_36_port, a(35) => 
                           final_first_level_0_35_port, a(34) => 
                           final_first_level_0_34_port, a(33) => 
                           final_first_level_0_33_port, a(32) => 
                           final_first_level_0_32_port, a(31) => 
                           final_first_level_0_31_port, a(30) => 
                           final_first_level_0_30_port, a(29) => 
                           final_first_level_0_29_port, a(28) => 
                           final_first_level_0_28_port, a(27) => 
                           final_first_level_0_27_port, a(26) => 
                           final_first_level_0_26_port, a(25) => 
                           final_first_level_0_25_port, a(24) => 
                           final_first_level_0_24_port, a(23) => 
                           final_first_level_0_23_port, a(22) => 
                           final_first_level_0_22_port, a(21) => 
                           final_first_level_0_21_port, a(20) => 
                           final_first_level_0_20_port, a(19) => 
                           final_first_level_0_19_port, a(18) => 
                           final_first_level_0_18_port, a(17) => 
                           final_first_level_0_17_port, a(16) => 
                           final_first_level_0_16_port, a(15) => 
                           final_first_level_0_15_port, a(14) => 
                           final_first_level_0_14_port, a(13) => 
                           final_first_level_0_13_port, a(12) => 
                           final_first_level_0_12_port, a(11) => 
                           final_first_level_0_11_port, a(10) => 
                           final_first_level_0_10_port, a(9) => 
                           final_first_level_0_9_port, a(8) => 
                           final_first_level_0_8_port, a(7) => 
                           final_first_level_0_7_port, a(6) => 
                           final_first_level_0_6_port, a(5) => 
                           final_first_level_0_5_port, a(4) => 
                           final_first_level_0_4_port, a(3) => 
                           final_first_level_0_3_port, a(2) => 
                           final_first_level_0_2_port, a(1) => 
                           final_first_level_0_1_port, a(0) => 
                           final_first_level_0_0_port, b(39) => 
                           final_first_level_1_39_port, b(38) => 
                           final_first_level_1_38_port, b(37) => 
                           final_first_level_1_37_port, b(36) => 
                           final_first_level_1_36_port, b(35) => 
                           final_first_level_1_35_port, b(34) => 
                           final_first_level_1_34_port, b(33) => 
                           final_first_level_1_33_port, b(32) => 
                           final_first_level_1_32_port, b(31) => 
                           final_first_level_1_31_port, b(30) => 
                           final_first_level_1_30_port, b(29) => 
                           final_first_level_1_29_port, b(28) => 
                           final_first_level_1_28_port, b(27) => 
                           final_first_level_1_27_port, b(26) => 
                           final_first_level_1_26_port, b(25) => 
                           final_first_level_1_25_port, b(24) => 
                           final_first_level_1_24_port, b(23) => 
                           final_first_level_1_23_port, b(22) => 
                           final_first_level_1_22_port, b(21) => 
                           final_first_level_1_21_port, b(20) => 
                           final_first_level_1_20_port, b(19) => 
                           final_first_level_1_19_port, b(18) => 
                           final_first_level_1_18_port, b(17) => 
                           final_first_level_1_17_port, b(16) => 
                           final_first_level_1_16_port, b(15) => 
                           final_first_level_1_15_port, b(14) => 
                           final_first_level_1_14_port, b(13) => 
                           final_first_level_1_13_port, b(12) => 
                           final_first_level_1_12_port, b(11) => 
                           final_first_level_1_11_port, b(10) => 
                           final_first_level_1_10_port, b(9) => 
                           final_first_level_1_9_port, b(8) => 
                           final_first_level_1_8_port, b(7) => 
                           final_first_level_1_7_port, b(6) => 
                           final_first_level_1_6_port, b(5) => 
                           final_first_level_1_5_port, b(4) => 
                           final_first_level_1_4_port, b(3) => 
                           final_first_level_1_3_port, b(2) => 
                           final_first_level_1_2_port, b(1) => 
                           final_first_level_1_1_port, b(0) => 
                           final_first_level_1_0_port, c(39) => 
                           final_first_level_2_39_port, c(38) => 
                           final_first_level_2_38_port, c(37) => 
                           final_first_level_2_37_port, c(36) => 
                           final_first_level_2_36_port, c(35) => 
                           final_first_level_2_35_port, c(34) => 
                           final_first_level_2_34_port, c(33) => 
                           final_first_level_2_33_port, c(32) => 
                           final_first_level_2_32_port, c(31) => 
                           final_first_level_2_31_port, c(30) => 
                           final_first_level_2_30_port, c(29) => 
                           final_first_level_2_29_port, c(28) => 
                           final_first_level_2_28_port, c(27) => 
                           final_first_level_2_27_port, c(26) => 
                           final_first_level_2_26_port, c(25) => 
                           final_first_level_2_25_port, c(24) => 
                           final_first_level_2_24_port, c(23) => 
                           final_first_level_2_23_port, c(22) => 
                           final_first_level_2_22_port, c(21) => 
                           final_first_level_2_21_port, c(20) => 
                           final_first_level_2_20_port, c(19) => 
                           final_first_level_2_19_port, c(18) => 
                           final_first_level_2_18_port, c(17) => 
                           final_first_level_2_17_port, c(16) => 
                           final_first_level_2_16_port, c(15) => 
                           final_first_level_2_15_port, c(14) => 
                           final_first_level_2_14_port, c(13) => 
                           final_first_level_2_13_port, c(12) => 
                           final_first_level_2_12_port, c(11) => 
                           final_first_level_2_11_port, c(10) => 
                           final_first_level_2_10_port, c(9) => 
                           final_first_level_2_9_port, c(8) => 
                           final_first_level_2_8_port, c(7) => 
                           final_first_level_2_7_port, c(6) => 
                           final_first_level_2_6_port, c(5) => 
                           final_first_level_2_5_port, c(4) => 
                           final_first_level_2_4_port, c(3) => 
                           final_first_level_2_3_port, c(2) => 
                           final_first_level_2_2_port, c(1) => 
                           final_first_level_2_1_port, c(0) => 
                           final_first_level_2_0_port, d(39) => 
                           final_first_level_3_39_port, d(38) => 
                           final_first_level_3_38_port, d(37) => 
                           final_first_level_3_37_port, d(36) => 
                           final_first_level_3_36_port, d(35) => 
                           final_first_level_3_35_port, d(34) => 
                           final_first_level_3_34_port, d(33) => 
                           final_first_level_3_33_port, d(32) => 
                           final_first_level_3_32_port, d(31) => 
                           final_first_level_3_31_port, d(30) => 
                           final_first_level_3_30_port, d(29) => 
                           final_first_level_3_29_port, d(28) => 
                           final_first_level_3_28_port, d(27) => 
                           final_first_level_3_27_port, d(26) => 
                           final_first_level_3_26_port, d(25) => 
                           final_first_level_3_25_port, d(24) => 
                           final_first_level_3_24_port, d(23) => 
                           final_first_level_3_23_port, d(22) => 
                           final_first_level_3_22_port, d(21) => 
                           final_first_level_3_21_port, d(20) => 
                           final_first_level_3_20_port, d(19) => 
                           final_first_level_3_19_port, d(18) => 
                           final_first_level_3_18_port, d(17) => 
                           final_first_level_3_17_port, d(16) => 
                           final_first_level_3_16_port, d(15) => 
                           final_first_level_3_15_port, d(14) => 
                           final_first_level_3_14_port, d(13) => 
                           final_first_level_3_13_port, d(12) => 
                           final_first_level_3_12_port, d(11) => 
                           final_first_level_3_11_port, d(10) => 
                           final_first_level_3_10_port, d(9) => 
                           final_first_level_3_9_port, d(8) => 
                           final_first_level_3_8_port, d(7) => 
                           final_first_level_3_7_port, d(6) => 
                           final_first_level_3_6_port, d(5) => 
                           final_first_level_3_5_port, d(4) => 
                           final_first_level_3_4_port, d(3) => 
                           final_first_level_3_3_port, d(2) => 
                           final_first_level_3_2_port, d(1) => 
                           final_first_level_3_1_port, d(0) => 
                           final_first_level_3_0_port, sel(1) => r2(4), sel(0) 
                           => r2(3), y(39) => n_1163, y(38) => 
                           final_first_level_mask_38_port, y(37) => 
                           final_first_level_mask_37_port, y(36) => 
                           final_first_level_mask_36_port, y(35) => 
                           final_first_level_mask_35_port, y(34) => 
                           final_first_level_mask_34_port, y(33) => 
                           final_first_level_mask_33_port, y(32) => 
                           final_first_level_mask_32_port, y(31) => 
                           final_first_level_mask_31_port, y(30) => 
                           final_first_level_mask_30_port, y(29) => 
                           final_first_level_mask_29_port, y(28) => 
                           final_first_level_mask_28_port, y(27) => 
                           final_first_level_mask_27_port, y(26) => 
                           final_first_level_mask_26_port, y(25) => 
                           final_first_level_mask_25_port, y(24) => 
                           final_first_level_mask_24_port, y(23) => 
                           final_first_level_mask_23_port, y(22) => 
                           final_first_level_mask_22_port, y(21) => 
                           final_first_level_mask_21_port, y(20) => 
                           final_first_level_mask_20_port, y(19) => 
                           final_first_level_mask_19_port, y(18) => 
                           final_first_level_mask_18_port, y(17) => 
                           final_first_level_mask_17_port, y(16) => 
                           final_first_level_mask_16_port, y(15) => 
                           final_first_level_mask_15_port, y(14) => 
                           final_first_level_mask_14_port, y(13) => 
                           final_first_level_mask_13_port, y(12) => 
                           final_first_level_mask_12_port, y(11) => 
                           final_first_level_mask_11_port, y(10) => 
                           final_first_level_mask_10_port, y(9) => 
                           final_first_level_mask_9_port, y(8) => 
                           final_first_level_mask_8_port, y(7) => 
                           final_first_level_mask_7_port, y(6) => 
                           final_first_level_mask_6_port, y(5) => 
                           final_first_level_mask_5_port, y(4) => 
                           final_first_level_mask_4_port, y(3) => 
                           final_first_level_mask_3_port, y(2) => 
                           final_first_level_mask_2_port, y(1) => 
                           final_first_level_mask_1_port, y(0) => 
                           final_first_level_mask_0_port);
   MUX81_level_3 : MUX81_N32 port map( a(31) => final_first_level_mask_31_port,
                           a(30) => final_first_level_mask_30_port, a(29) => 
                           final_first_level_mask_29_port, a(28) => 
                           final_first_level_mask_28_port, a(27) => 
                           final_first_level_mask_27_port, a(26) => 
                           final_first_level_mask_26_port, a(25) => 
                           final_first_level_mask_25_port, a(24) => 
                           final_first_level_mask_24_port, a(23) => 
                           final_first_level_mask_23_port, a(22) => 
                           final_first_level_mask_22_port, a(21) => 
                           final_first_level_mask_21_port, a(20) => 
                           final_first_level_mask_20_port, a(19) => 
                           final_first_level_mask_19_port, a(18) => 
                           final_first_level_mask_18_port, a(17) => 
                           final_first_level_mask_17_port, a(16) => 
                           final_first_level_mask_16_port, a(15) => 
                           final_first_level_mask_15_port, a(14) => 
                           final_first_level_mask_14_port, a(13) => 
                           final_first_level_mask_13_port, a(12) => 
                           final_first_level_mask_12_port, a(11) => 
                           final_first_level_mask_11_port, a(10) => 
                           final_first_level_mask_10_port, a(9) => 
                           final_first_level_mask_9_port, a(8) => 
                           final_first_level_mask_8_port, a(7) => 
                           final_first_level_mask_7_port, a(6) => 
                           final_first_level_mask_6_port, a(5) => 
                           final_first_level_mask_5_port, a(4) => 
                           final_first_level_mask_4_port, a(3) => 
                           final_first_level_mask_3_port, a(2) => 
                           final_first_level_mask_2_port, a(1) => 
                           final_first_level_mask_1_port, a(0) => 
                           final_first_level_mask_0_port, b(31) => 
                           final_first_level_mask_32_port, b(30) => 
                           final_first_level_mask_31_port, b(29) => 
                           final_first_level_mask_30_port, b(28) => 
                           final_first_level_mask_29_port, b(27) => 
                           final_first_level_mask_28_port, b(26) => 
                           final_first_level_mask_27_port, b(25) => 
                           final_first_level_mask_26_port, b(24) => 
                           final_first_level_mask_25_port, b(23) => 
                           final_first_level_mask_24_port, b(22) => 
                           final_first_level_mask_23_port, b(21) => 
                           final_first_level_mask_22_port, b(20) => 
                           final_first_level_mask_21_port, b(19) => 
                           final_first_level_mask_20_port, b(18) => 
                           final_first_level_mask_19_port, b(17) => 
                           final_first_level_mask_18_port, b(16) => 
                           final_first_level_mask_17_port, b(15) => 
                           final_first_level_mask_16_port, b(14) => 
                           final_first_level_mask_15_port, b(13) => 
                           final_first_level_mask_14_port, b(12) => 
                           final_first_level_mask_13_port, b(11) => 
                           final_first_level_mask_12_port, b(10) => 
                           final_first_level_mask_11_port, b(9) => 
                           final_first_level_mask_10_port, b(8) => 
                           final_first_level_mask_9_port, b(7) => 
                           final_first_level_mask_8_port, b(6) => 
                           final_first_level_mask_7_port, b(5) => 
                           final_first_level_mask_6_port, b(4) => 
                           final_first_level_mask_5_port, b(3) => 
                           final_first_level_mask_4_port, b(2) => 
                           final_first_level_mask_3_port, b(1) => 
                           final_first_level_mask_2_port, b(0) => 
                           final_first_level_mask_1_port, c(31) => 
                           final_first_level_mask_33_port, c(30) => 
                           final_first_level_mask_32_port, c(29) => 
                           final_first_level_mask_31_port, c(28) => 
                           final_first_level_mask_30_port, c(27) => 
                           final_first_level_mask_29_port, c(26) => 
                           final_first_level_mask_28_port, c(25) => 
                           final_first_level_mask_27_port, c(24) => 
                           final_first_level_mask_26_port, c(23) => 
                           final_first_level_mask_25_port, c(22) => 
                           final_first_level_mask_24_port, c(21) => 
                           final_first_level_mask_23_port, c(20) => 
                           final_first_level_mask_22_port, c(19) => 
                           final_first_level_mask_21_port, c(18) => 
                           final_first_level_mask_20_port, c(17) => 
                           final_first_level_mask_19_port, c(16) => 
                           final_first_level_mask_18_port, c(15) => 
                           final_first_level_mask_17_port, c(14) => 
                           final_first_level_mask_16_port, c(13) => 
                           final_first_level_mask_15_port, c(12) => 
                           final_first_level_mask_14_port, c(11) => 
                           final_first_level_mask_13_port, c(10) => 
                           final_first_level_mask_12_port, c(9) => 
                           final_first_level_mask_11_port, c(8) => 
                           final_first_level_mask_10_port, c(7) => 
                           final_first_level_mask_9_port, c(6) => 
                           final_first_level_mask_8_port, c(5) => 
                           final_first_level_mask_7_port, c(4) => 
                           final_first_level_mask_6_port, c(3) => 
                           final_first_level_mask_5_port, c(2) => 
                           final_first_level_mask_4_port, c(1) => 
                           final_first_level_mask_3_port, c(0) => 
                           final_first_level_mask_2_port, d(31) => 
                           final_first_level_mask_34_port, d(30) => 
                           final_first_level_mask_33_port, d(29) => 
                           final_first_level_mask_32_port, d(28) => 
                           final_first_level_mask_31_port, d(27) => 
                           final_first_level_mask_30_port, d(26) => 
                           final_first_level_mask_29_port, d(25) => 
                           final_first_level_mask_28_port, d(24) => 
                           final_first_level_mask_27_port, d(23) => 
                           final_first_level_mask_26_port, d(22) => 
                           final_first_level_mask_25_port, d(21) => 
                           final_first_level_mask_24_port, d(20) => 
                           final_first_level_mask_23_port, d(19) => 
                           final_first_level_mask_22_port, d(18) => 
                           final_first_level_mask_21_port, d(17) => 
                           final_first_level_mask_20_port, d(16) => 
                           final_first_level_mask_19_port, d(15) => 
                           final_first_level_mask_18_port, d(14) => 
                           final_first_level_mask_17_port, d(13) => 
                           final_first_level_mask_16_port, d(12) => 
                           final_first_level_mask_15_port, d(11) => 
                           final_first_level_mask_14_port, d(10) => 
                           final_first_level_mask_13_port, d(9) => 
                           final_first_level_mask_12_port, d(8) => 
                           final_first_level_mask_11_port, d(7) => 
                           final_first_level_mask_10_port, d(6) => 
                           final_first_level_mask_9_port, d(5) => 
                           final_first_level_mask_8_port, d(4) => 
                           final_first_level_mask_7_port, d(3) => 
                           final_first_level_mask_6_port, d(2) => 
                           final_first_level_mask_5_port, d(1) => 
                           final_first_level_mask_4_port, d(0) => 
                           final_first_level_mask_3_port, e(31) => 
                           final_first_level_mask_35_port, e(30) => 
                           final_first_level_mask_34_port, e(29) => 
                           final_first_level_mask_33_port, e(28) => 
                           final_first_level_mask_32_port, e(27) => 
                           final_first_level_mask_31_port, e(26) => 
                           final_first_level_mask_30_port, e(25) => 
                           final_first_level_mask_29_port, e(24) => 
                           final_first_level_mask_28_port, e(23) => 
                           final_first_level_mask_27_port, e(22) => 
                           final_first_level_mask_26_port, e(21) => 
                           final_first_level_mask_25_port, e(20) => 
                           final_first_level_mask_24_port, e(19) => 
                           final_first_level_mask_23_port, e(18) => 
                           final_first_level_mask_22_port, e(17) => 
                           final_first_level_mask_21_port, e(16) => 
                           final_first_level_mask_20_port, e(15) => 
                           final_first_level_mask_19_port, e(14) => 
                           final_first_level_mask_18_port, e(13) => 
                           final_first_level_mask_17_port, e(12) => 
                           final_first_level_mask_16_port, e(11) => 
                           final_first_level_mask_15_port, e(10) => 
                           final_first_level_mask_14_port, e(9) => 
                           final_first_level_mask_13_port, e(8) => 
                           final_first_level_mask_12_port, e(7) => 
                           final_first_level_mask_11_port, e(6) => 
                           final_first_level_mask_10_port, e(5) => 
                           final_first_level_mask_9_port, e(4) => 
                           final_first_level_mask_8_port, e(3) => 
                           final_first_level_mask_7_port, e(2) => 
                           final_first_level_mask_6_port, e(1) => 
                           final_first_level_mask_5_port, e(0) => 
                           final_first_level_mask_4_port, f(31) => 
                           final_first_level_mask_36_port, f(30) => 
                           final_first_level_mask_35_port, f(29) => 
                           final_first_level_mask_34_port, f(28) => 
                           final_first_level_mask_33_port, f(27) => 
                           final_first_level_mask_32_port, f(26) => 
                           final_first_level_mask_31_port, f(25) => 
                           final_first_level_mask_30_port, f(24) => 
                           final_first_level_mask_29_port, f(23) => 
                           final_first_level_mask_28_port, f(22) => 
                           final_first_level_mask_27_port, f(21) => 
                           final_first_level_mask_26_port, f(20) => 
                           final_first_level_mask_25_port, f(19) => 
                           final_first_level_mask_24_port, f(18) => 
                           final_first_level_mask_23_port, f(17) => 
                           final_first_level_mask_22_port, f(16) => 
                           final_first_level_mask_21_port, f(15) => 
                           final_first_level_mask_20_port, f(14) => 
                           final_first_level_mask_19_port, f(13) => 
                           final_first_level_mask_18_port, f(12) => 
                           final_first_level_mask_17_port, f(11) => 
                           final_first_level_mask_16_port, f(10) => 
                           final_first_level_mask_15_port, f(9) => 
                           final_first_level_mask_14_port, f(8) => 
                           final_first_level_mask_13_port, f(7) => 
                           final_first_level_mask_12_port, f(6) => 
                           final_first_level_mask_11_port, f(5) => 
                           final_first_level_mask_10_port, f(4) => 
                           final_first_level_mask_9_port, f(3) => 
                           final_first_level_mask_8_port, f(2) => 
                           final_first_level_mask_7_port, f(1) => 
                           final_first_level_mask_6_port, f(0) => 
                           final_first_level_mask_5_port, g(31) => 
                           final_first_level_mask_37_port, g(30) => 
                           final_first_level_mask_36_port, g(29) => 
                           final_first_level_mask_35_port, g(28) => 
                           final_first_level_mask_34_port, g(27) => 
                           final_first_level_mask_33_port, g(26) => 
                           final_first_level_mask_32_port, g(25) => 
                           final_first_level_mask_31_port, g(24) => 
                           final_first_level_mask_30_port, g(23) => 
                           final_first_level_mask_29_port, g(22) => 
                           final_first_level_mask_28_port, g(21) => 
                           final_first_level_mask_27_port, g(20) => 
                           final_first_level_mask_26_port, g(19) => 
                           final_first_level_mask_25_port, g(18) => 
                           final_first_level_mask_24_port, g(17) => 
                           final_first_level_mask_23_port, g(16) => 
                           final_first_level_mask_22_port, g(15) => 
                           final_first_level_mask_21_port, g(14) => 
                           final_first_level_mask_20_port, g(13) => 
                           final_first_level_mask_19_port, g(12) => 
                           final_first_level_mask_18_port, g(11) => 
                           final_first_level_mask_17_port, g(10) => 
                           final_first_level_mask_16_port, g(9) => 
                           final_first_level_mask_15_port, g(8) => 
                           final_first_level_mask_14_port, g(7) => 
                           final_first_level_mask_13_port, g(6) => 
                           final_first_level_mask_12_port, g(5) => 
                           final_first_level_mask_11_port, g(4) => 
                           final_first_level_mask_10_port, g(3) => 
                           final_first_level_mask_9_port, g(2) => 
                           final_first_level_mask_8_port, g(1) => 
                           final_first_level_mask_7_port, g(0) => 
                           final_first_level_mask_6_port, h(31) => 
                           final_first_level_mask_38_port, h(30) => 
                           final_first_level_mask_37_port, h(29) => 
                           final_first_level_mask_36_port, h(28) => 
                           final_first_level_mask_35_port, h(27) => 
                           final_first_level_mask_34_port, h(26) => 
                           final_first_level_mask_33_port, h(25) => 
                           final_first_level_mask_32_port, h(24) => 
                           final_first_level_mask_31_port, h(23) => 
                           final_first_level_mask_30_port, h(22) => 
                           final_first_level_mask_29_port, h(21) => 
                           final_first_level_mask_28_port, h(20) => 
                           final_first_level_mask_27_port, h(19) => 
                           final_first_level_mask_26_port, h(18) => 
                           final_first_level_mask_25_port, h(17) => 
                           final_first_level_mask_24_port, h(16) => 
                           final_first_level_mask_23_port, h(15) => 
                           final_first_level_mask_22_port, h(14) => 
                           final_first_level_mask_21_port, h(13) => 
                           final_first_level_mask_20_port, h(12) => 
                           final_first_level_mask_19_port, h(11) => 
                           final_first_level_mask_18_port, h(10) => 
                           final_first_level_mask_17_port, h(9) => 
                           final_first_level_mask_16_port, h(8) => 
                           final_first_level_mask_15_port, h(7) => 
                           final_first_level_mask_14_port, h(6) => 
                           final_first_level_mask_13_port, h(5) => 
                           final_first_level_mask_12_port, h(4) => 
                           final_first_level_mask_11_port, h(3) => 
                           final_first_level_mask_10_port, h(2) => 
                           final_first_level_mask_9_port, h(1) => 
                           final_first_level_mask_8_port, h(0) => 
                           final_first_level_mask_7_port, sel(2) => 
                           third_level_sel_2_port, sel(1) => 
                           third_level_sel_1_port, sel(0) => 
                           third_level_sel_0_port, y(31) => shifted_out(31), 
                           y(30) => shifted_out(30), y(29) => shifted_out(29), 
                           y(28) => shifted_out(28), y(27) => shifted_out(27), 
                           y(26) => shifted_out(26), y(25) => shifted_out(25), 
                           y(24) => shifted_out(24), y(23) => shifted_out(23), 
                           y(22) => shifted_out(22), y(21) => shifted_out(21), 
                           y(20) => shifted_out(20), y(19) => shifted_out(19), 
                           y(18) => shifted_out(18), y(17) => shifted_out(17), 
                           y(16) => shifted_out(16), y(15) => shifted_out(15), 
                           y(14) => shifted_out(14), y(13) => shifted_out(13), 
                           y(12) => shifted_out(12), y(11) => shifted_out(11), 
                           y(10) => shifted_out(10), y(9) => shifted_out(9), 
                           y(8) => shifted_out(8), y(7) => shifted_out(7), y(6)
                           => shifted_out(6), y(5) => shifted_out(5), y(4) => 
                           shifted_out(4), y(3) => shifted_out(3), y(2) => 
                           shifted_out(2), y(1) => shifted_out(1), y(0) => 
                           shifted_out(0));
   U2 : AND2_X4 port map( A1 => r1(31), A2 => conf(1), ZN => 
                           right_first_level_3_39_port);
   U3 : XOR2_X1 port map( A => r2(2), B => conf(0), Z => third_level_sel_2_port
                           );
   U4 : XOR2_X1 port map( A => r2(1), B => conf(0), Z => third_level_sel_1_port
                           );
   U5 : XOR2_X1 port map( A => r2(0), B => conf(0), Z => third_level_sel_0_port
                           );

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity boothmul_NBIT32_N16_M16 is

   port( a, b : in std_logic_vector (15 downto 0);  mul : out std_logic_vector 
         (31 downto 0));

end boothmul_NBIT32_N16_M16;

architecture SYN_structural of boothmul_NBIT32_N16_M16 is

   component rca_signed_NBIT32_1
      port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_1
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT7
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   component rca_signed_NBIT32_2
      port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_2
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT6
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   component rca_signed_NBIT32_3
      port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_3
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT5
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   component rca_signed_NBIT32_4
      port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_4
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT4
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   component rca_signed_NBIT32_5
      port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_5
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT3
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   component rca_signed_NBIT32_6
      port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_6
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT2
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   component rca_signed_NBIT32_0
      port( a, b : in std_logic_vector (31 downto 0);  c : out std_logic;  s : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_7
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT1
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   component vp_NBIT32_0
      port( pos_a, neg_a, pos_2a, neg_2a : in std_logic_vector (31 downto 0);  
            sel : in std_logic_vector (2 downto 0);  s_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_NBIT32_SHIFT0
      port( a : in std_logic_vector (15 downto 0);  pos_a, neg_a, pos_2a, 
            neg_2a : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, neg_2av_7_31_port, neg_2av_7_30_port, 
      neg_2av_7_29_port, neg_2av_7_28_port, neg_2av_7_27_port, 
      neg_2av_7_26_port, neg_2av_7_25_port, neg_2av_7_24_port, 
      neg_2av_7_23_port, neg_2av_7_22_port, neg_2av_7_21_port, 
      neg_2av_7_20_port, neg_2av_7_19_port, neg_2av_7_18_port, 
      neg_2av_7_17_port, neg_2av_7_16_port, neg_2av_7_15_port, 
      neg_2av_7_14_port, neg_2av_7_13_port, neg_2av_7_12_port, 
      neg_2av_7_11_port, neg_2av_7_10_port, neg_2av_7_9_port, neg_2av_7_8_port,
      neg_2av_7_7_port, neg_2av_7_6_port, neg_2av_7_5_port, neg_2av_7_4_port, 
      neg_2av_7_3_port, neg_2av_7_2_port, neg_2av_7_1_port, neg_2av_7_0_port, 
      neg_2av_6_31_port, neg_2av_6_30_port, neg_2av_6_29_port, 
      neg_2av_6_28_port, neg_2av_6_27_port, neg_2av_6_26_port, 
      neg_2av_6_25_port, neg_2av_6_24_port, neg_2av_6_23_port, 
      neg_2av_6_22_port, neg_2av_6_21_port, neg_2av_6_20_port, 
      neg_2av_6_19_port, neg_2av_6_18_port, neg_2av_6_17_port, 
      neg_2av_6_16_port, neg_2av_6_15_port, neg_2av_6_14_port, 
      neg_2av_6_13_port, neg_2av_6_12_port, neg_2av_6_11_port, 
      neg_2av_6_10_port, neg_2av_6_9_port, neg_2av_6_8_port, neg_2av_6_7_port, 
      neg_2av_6_6_port, neg_2av_6_5_port, neg_2av_6_4_port, neg_2av_6_3_port, 
      neg_2av_6_2_port, neg_2av_6_1_port, neg_2av_6_0_port, neg_2av_5_31_port, 
      neg_2av_5_30_port, neg_2av_5_29_port, neg_2av_5_28_port, 
      neg_2av_5_27_port, neg_2av_5_26_port, neg_2av_5_25_port, 
      neg_2av_5_24_port, neg_2av_5_23_port, neg_2av_5_22_port, 
      neg_2av_5_21_port, neg_2av_5_20_port, neg_2av_5_19_port, 
      neg_2av_5_18_port, neg_2av_5_17_port, neg_2av_5_16_port, 
      neg_2av_5_15_port, neg_2av_5_14_port, neg_2av_5_13_port, 
      neg_2av_5_12_port, neg_2av_5_11_port, neg_2av_5_10_port, neg_2av_5_9_port
      , neg_2av_5_8_port, neg_2av_5_7_port, neg_2av_5_6_port, neg_2av_5_5_port,
      neg_2av_5_4_port, neg_2av_5_3_port, neg_2av_5_2_port, neg_2av_5_1_port, 
      neg_2av_5_0_port, neg_2av_4_31_port, neg_2av_4_30_port, neg_2av_4_29_port
      , neg_2av_4_28_port, neg_2av_4_27_port, neg_2av_4_26_port, 
      neg_2av_4_25_port, neg_2av_4_24_port, neg_2av_4_23_port, 
      neg_2av_4_22_port, neg_2av_4_21_port, neg_2av_4_20_port, 
      neg_2av_4_19_port, neg_2av_4_18_port, neg_2av_4_17_port, 
      neg_2av_4_16_port, neg_2av_4_15_port, neg_2av_4_14_port, 
      neg_2av_4_13_port, neg_2av_4_12_port, neg_2av_4_11_port, 
      neg_2av_4_10_port, neg_2av_4_9_port, neg_2av_4_8_port, neg_2av_4_7_port, 
      neg_2av_4_6_port, neg_2av_4_5_port, neg_2av_4_4_port, neg_2av_4_3_port, 
      neg_2av_4_2_port, neg_2av_4_1_port, neg_2av_4_0_port, neg_2av_3_31_port, 
      neg_2av_3_30_port, neg_2av_3_29_port, neg_2av_3_28_port, 
      neg_2av_3_27_port, neg_2av_3_26_port, neg_2av_3_25_port, 
      neg_2av_3_24_port, neg_2av_3_23_port, neg_2av_3_22_port, 
      neg_2av_3_21_port, neg_2av_3_20_port, neg_2av_3_19_port, 
      neg_2av_3_18_port, neg_2av_3_17_port, neg_2av_3_16_port, 
      neg_2av_3_15_port, neg_2av_3_14_port, neg_2av_3_13_port, 
      neg_2av_3_12_port, neg_2av_3_11_port, neg_2av_3_10_port, neg_2av_3_9_port
      , neg_2av_3_8_port, neg_2av_3_7_port, neg_2av_3_6_port, neg_2av_3_5_port,
      neg_2av_3_4_port, neg_2av_3_3_port, neg_2av_3_2_port, neg_2av_3_1_port, 
      neg_2av_3_0_port, neg_2av_2_31_port, neg_2av_2_30_port, neg_2av_2_29_port
      , neg_2av_2_28_port, neg_2av_2_27_port, neg_2av_2_26_port, 
      neg_2av_2_25_port, neg_2av_2_24_port, neg_2av_2_23_port, 
      neg_2av_2_22_port, neg_2av_2_21_port, neg_2av_2_20_port, 
      neg_2av_2_19_port, neg_2av_2_18_port, neg_2av_2_17_port, 
      neg_2av_2_16_port, neg_2av_2_15_port, neg_2av_2_14_port, 
      neg_2av_2_13_port, neg_2av_2_12_port, neg_2av_2_11_port, 
      neg_2av_2_10_port, neg_2av_2_9_port, neg_2av_2_8_port, neg_2av_2_7_port, 
      neg_2av_2_6_port, neg_2av_2_5_port, neg_2av_2_4_port, neg_2av_2_3_port, 
      neg_2av_2_2_port, neg_2av_2_1_port, neg_2av_2_0_port, neg_2av_1_31_port, 
      neg_2av_1_30_port, neg_2av_1_29_port, neg_2av_1_28_port, 
      neg_2av_1_27_port, neg_2av_1_26_port, neg_2av_1_25_port, 
      neg_2av_1_24_port, neg_2av_1_23_port, neg_2av_1_22_port, 
      neg_2av_1_21_port, neg_2av_1_20_port, neg_2av_1_19_port, 
      neg_2av_1_18_port, neg_2av_1_17_port, neg_2av_1_16_port, 
      neg_2av_1_15_port, neg_2av_1_14_port, neg_2av_1_13_port, 
      neg_2av_1_12_port, neg_2av_1_11_port, neg_2av_1_10_port, neg_2av_1_9_port
      , neg_2av_1_8_port, neg_2av_1_7_port, neg_2av_1_6_port, neg_2av_1_5_port,
      neg_2av_1_4_port, neg_2av_1_3_port, neg_2av_1_2_port, neg_2av_1_1_port, 
      neg_2av_1_0_port, neg_2av_0_31_port, neg_2av_0_30_port, neg_2av_0_29_port
      , neg_2av_0_28_port, neg_2av_0_27_port, neg_2av_0_26_port, 
      neg_2av_0_25_port, neg_2av_0_24_port, neg_2av_0_23_port, 
      neg_2av_0_22_port, neg_2av_0_21_port, neg_2av_0_20_port, 
      neg_2av_0_19_port, neg_2av_0_18_port, neg_2av_0_17_port, 
      neg_2av_0_16_port, neg_2av_0_15_port, neg_2av_0_14_port, 
      neg_2av_0_13_port, neg_2av_0_12_port, neg_2av_0_11_port, 
      neg_2av_0_10_port, neg_2av_0_9_port, neg_2av_0_8_port, neg_2av_0_7_port, 
      neg_2av_0_6_port, neg_2av_0_5_port, neg_2av_0_4_port, neg_2av_0_3_port, 
      neg_2av_0_2_port, neg_2av_0_1_port, neg_2av_0_0_port, pos_2av_7_31_port, 
      pos_2av_7_30_port, pos_2av_7_29_port, pos_2av_7_28_port, 
      pos_2av_7_27_port, pos_2av_7_26_port, pos_2av_7_25_port, 
      pos_2av_7_24_port, pos_2av_7_23_port, pos_2av_7_22_port, 
      pos_2av_7_21_port, pos_2av_7_20_port, pos_2av_7_19_port, 
      pos_2av_7_18_port, pos_2av_7_17_port, pos_2av_7_16_port, 
      pos_2av_7_15_port, pos_2av_7_14_port, pos_2av_7_13_port, 
      pos_2av_7_12_port, pos_2av_7_11_port, pos_2av_7_10_port, pos_2av_7_9_port
      , pos_2av_7_8_port, pos_2av_7_7_port, pos_2av_7_6_port, pos_2av_7_5_port,
      pos_2av_7_4_port, pos_2av_7_3_port, pos_2av_7_2_port, pos_2av_7_1_port, 
      pos_2av_7_0_port, pos_2av_6_31_port, pos_2av_6_30_port, pos_2av_6_29_port
      , pos_2av_6_28_port, pos_2av_6_27_port, pos_2av_6_26_port, 
      pos_2av_6_25_port, pos_2av_6_24_port, pos_2av_6_23_port, 
      pos_2av_6_22_port, pos_2av_6_21_port, pos_2av_6_20_port, 
      pos_2av_6_19_port, pos_2av_6_18_port, pos_2av_6_17_port, 
      pos_2av_6_16_port, pos_2av_6_15_port, pos_2av_6_14_port, 
      pos_2av_6_13_port, pos_2av_6_12_port, pos_2av_6_11_port, 
      pos_2av_6_10_port, pos_2av_6_9_port, pos_2av_6_8_port, pos_2av_6_7_port, 
      pos_2av_6_6_port, pos_2av_6_5_port, pos_2av_6_4_port, pos_2av_6_3_port, 
      pos_2av_6_2_port, pos_2av_6_1_port, pos_2av_6_0_port, pos_2av_5_31_port, 
      pos_2av_5_30_port, pos_2av_5_29_port, pos_2av_5_28_port, 
      pos_2av_5_27_port, pos_2av_5_26_port, pos_2av_5_25_port, 
      pos_2av_5_24_port, pos_2av_5_23_port, pos_2av_5_22_port, 
      pos_2av_5_21_port, pos_2av_5_20_port, pos_2av_5_19_port, 
      pos_2av_5_18_port, pos_2av_5_17_port, pos_2av_5_16_port, 
      pos_2av_5_15_port, pos_2av_5_14_port, pos_2av_5_13_port, 
      pos_2av_5_12_port, pos_2av_5_11_port, pos_2av_5_10_port, pos_2av_5_9_port
      , pos_2av_5_8_port, pos_2av_5_7_port, pos_2av_5_6_port, pos_2av_5_5_port,
      pos_2av_5_4_port, pos_2av_5_3_port, pos_2av_5_2_port, pos_2av_5_1_port, 
      pos_2av_5_0_port, pos_2av_4_31_port, pos_2av_4_30_port, pos_2av_4_29_port
      , pos_2av_4_28_port, pos_2av_4_27_port, pos_2av_4_26_port, 
      pos_2av_4_25_port, pos_2av_4_24_port, pos_2av_4_23_port, 
      pos_2av_4_22_port, pos_2av_4_21_port, pos_2av_4_20_port, 
      pos_2av_4_19_port, pos_2av_4_18_port, pos_2av_4_17_port, 
      pos_2av_4_16_port, pos_2av_4_15_port, pos_2av_4_14_port, 
      pos_2av_4_13_port, pos_2av_4_12_port, pos_2av_4_11_port, 
      pos_2av_4_10_port, pos_2av_4_9_port, pos_2av_4_8_port, pos_2av_4_7_port, 
      pos_2av_4_6_port, pos_2av_4_5_port, pos_2av_4_4_port, pos_2av_4_3_port, 
      pos_2av_4_2_port, pos_2av_4_1_port, pos_2av_4_0_port, pos_2av_3_31_port, 
      pos_2av_3_30_port, pos_2av_3_29_port, pos_2av_3_28_port, 
      pos_2av_3_27_port, pos_2av_3_26_port, pos_2av_3_25_port, 
      pos_2av_3_24_port, pos_2av_3_23_port, pos_2av_3_22_port, 
      pos_2av_3_21_port, pos_2av_3_20_port, pos_2av_3_19_port, 
      pos_2av_3_18_port, pos_2av_3_17_port, pos_2av_3_16_port, 
      pos_2av_3_15_port, pos_2av_3_14_port, pos_2av_3_13_port, 
      pos_2av_3_12_port, pos_2av_3_11_port, pos_2av_3_10_port, pos_2av_3_9_port
      , pos_2av_3_8_port, pos_2av_3_7_port, pos_2av_3_6_port, pos_2av_3_5_port,
      pos_2av_3_4_port, pos_2av_3_3_port, pos_2av_3_2_port, pos_2av_3_1_port, 
      pos_2av_3_0_port, pos_2av_2_31_port, pos_2av_2_30_port, pos_2av_2_29_port
      , pos_2av_2_28_port, pos_2av_2_27_port, pos_2av_2_26_port, 
      pos_2av_2_25_port, pos_2av_2_24_port, pos_2av_2_23_port, 
      pos_2av_2_22_port, pos_2av_2_21_port, pos_2av_2_20_port, 
      pos_2av_2_19_port, pos_2av_2_18_port, pos_2av_2_17_port, 
      pos_2av_2_16_port, pos_2av_2_15_port, pos_2av_2_14_port, 
      pos_2av_2_13_port, pos_2av_2_12_port, pos_2av_2_11_port, 
      pos_2av_2_10_port, pos_2av_2_9_port, pos_2av_2_8_port, pos_2av_2_7_port, 
      pos_2av_2_6_port, pos_2av_2_5_port, pos_2av_2_4_port, pos_2av_2_3_port, 
      pos_2av_2_2_port, pos_2av_2_1_port, pos_2av_2_0_port, pos_2av_1_31_port, 
      pos_2av_1_30_port, pos_2av_1_29_port, pos_2av_1_28_port, 
      pos_2av_1_27_port, pos_2av_1_26_port, pos_2av_1_25_port, 
      pos_2av_1_24_port, pos_2av_1_23_port, pos_2av_1_22_port, 
      pos_2av_1_21_port, pos_2av_1_20_port, pos_2av_1_19_port, 
      pos_2av_1_18_port, pos_2av_1_17_port, pos_2av_1_16_port, 
      pos_2av_1_15_port, pos_2av_1_14_port, pos_2av_1_13_port, 
      pos_2av_1_12_port, pos_2av_1_11_port, pos_2av_1_10_port, pos_2av_1_9_port
      , pos_2av_1_8_port, pos_2av_1_7_port, pos_2av_1_6_port, pos_2av_1_5_port,
      pos_2av_1_4_port, pos_2av_1_3_port, pos_2av_1_2_port, pos_2av_1_1_port, 
      pos_2av_1_0_port, pos_2av_0_31_port, pos_2av_0_30_port, pos_2av_0_29_port
      , pos_2av_0_28_port, pos_2av_0_27_port, pos_2av_0_26_port, 
      pos_2av_0_25_port, pos_2av_0_24_port, pos_2av_0_23_port, 
      pos_2av_0_22_port, pos_2av_0_21_port, pos_2av_0_20_port, 
      pos_2av_0_19_port, pos_2av_0_18_port, pos_2av_0_17_port, 
      pos_2av_0_16_port, pos_2av_0_15_port, pos_2av_0_14_port, 
      pos_2av_0_13_port, pos_2av_0_12_port, pos_2av_0_11_port, 
      pos_2av_0_10_port, pos_2av_0_9_port, pos_2av_0_8_port, pos_2av_0_7_port, 
      pos_2av_0_6_port, pos_2av_0_5_port, pos_2av_0_4_port, pos_2av_0_3_port, 
      pos_2av_0_2_port, pos_2av_0_1_port, pos_2av_0_0_port, neg_av_7_31_port, 
      neg_av_7_30_port, neg_av_7_29_port, neg_av_7_28_port, neg_av_7_27_port, 
      neg_av_7_26_port, neg_av_7_25_port, neg_av_7_24_port, neg_av_7_23_port, 
      neg_av_7_22_port, neg_av_7_21_port, neg_av_7_20_port, neg_av_7_19_port, 
      neg_av_7_18_port, neg_av_7_17_port, neg_av_7_16_port, neg_av_7_15_port, 
      neg_av_7_14_port, neg_av_7_13_port, neg_av_7_12_port, neg_av_7_11_port, 
      neg_av_7_10_port, neg_av_7_9_port, neg_av_7_8_port, neg_av_7_7_port, 
      neg_av_7_6_port, neg_av_7_5_port, neg_av_7_4_port, neg_av_7_3_port, 
      neg_av_7_2_port, neg_av_7_1_port, neg_av_7_0_port, neg_av_6_31_port, 
      neg_av_6_30_port, neg_av_6_29_port, neg_av_6_28_port, neg_av_6_27_port, 
      neg_av_6_26_port, neg_av_6_25_port, neg_av_6_24_port, neg_av_6_23_port, 
      neg_av_6_22_port, neg_av_6_21_port, neg_av_6_20_port, neg_av_6_19_port, 
      neg_av_6_18_port, neg_av_6_17_port, neg_av_6_16_port, neg_av_6_15_port, 
      neg_av_6_14_port, neg_av_6_13_port, neg_av_6_12_port, neg_av_6_11_port, 
      neg_av_6_10_port, neg_av_6_9_port, neg_av_6_8_port, neg_av_6_7_port, 
      neg_av_6_6_port, neg_av_6_5_port, neg_av_6_4_port, neg_av_6_3_port, 
      neg_av_6_2_port, neg_av_6_1_port, neg_av_6_0_port, neg_av_5_31_port, 
      neg_av_5_30_port, neg_av_5_29_port, neg_av_5_28_port, neg_av_5_27_port, 
      neg_av_5_26_port, neg_av_5_25_port, neg_av_5_24_port, neg_av_5_23_port, 
      neg_av_5_22_port, neg_av_5_21_port, neg_av_5_20_port, neg_av_5_19_port, 
      neg_av_5_18_port, neg_av_5_17_port, neg_av_5_16_port, neg_av_5_15_port, 
      neg_av_5_14_port, neg_av_5_13_port, neg_av_5_12_port, neg_av_5_11_port, 
      neg_av_5_10_port, neg_av_5_9_port, neg_av_5_8_port, neg_av_5_7_port, 
      neg_av_5_6_port, neg_av_5_5_port, neg_av_5_4_port, neg_av_5_3_port, 
      neg_av_5_2_port, neg_av_5_1_port, neg_av_5_0_port, neg_av_4_31_port, 
      neg_av_4_30_port, neg_av_4_29_port, neg_av_4_28_port, neg_av_4_27_port, 
      neg_av_4_26_port, neg_av_4_25_port, neg_av_4_24_port, neg_av_4_23_port, 
      neg_av_4_22_port, neg_av_4_21_port, neg_av_4_20_port, neg_av_4_19_port, 
      neg_av_4_18_port, neg_av_4_17_port, neg_av_4_16_port, neg_av_4_15_port, 
      neg_av_4_14_port, neg_av_4_13_port, neg_av_4_12_port, neg_av_4_11_port, 
      neg_av_4_10_port, neg_av_4_9_port, neg_av_4_8_port, neg_av_4_7_port, 
      neg_av_4_6_port, neg_av_4_5_port, neg_av_4_4_port, neg_av_4_3_port, 
      neg_av_4_2_port, neg_av_4_1_port, neg_av_4_0_port, neg_av_3_31_port, 
      neg_av_3_30_port, neg_av_3_29_port, neg_av_3_28_port, neg_av_3_27_port, 
      neg_av_3_26_port, neg_av_3_25_port, neg_av_3_24_port, neg_av_3_23_port, 
      neg_av_3_22_port, neg_av_3_21_port, neg_av_3_20_port, neg_av_3_19_port, 
      neg_av_3_18_port, neg_av_3_17_port, neg_av_3_16_port, neg_av_3_15_port, 
      neg_av_3_14_port, neg_av_3_13_port, neg_av_3_12_port, neg_av_3_11_port, 
      neg_av_3_10_port, neg_av_3_9_port, neg_av_3_8_port, neg_av_3_7_port, 
      neg_av_3_6_port, neg_av_3_5_port, neg_av_3_4_port, neg_av_3_3_port, 
      neg_av_3_2_port, neg_av_3_1_port, neg_av_3_0_port, neg_av_2_31_port, 
      neg_av_2_30_port, neg_av_2_29_port, neg_av_2_28_port, neg_av_2_27_port, 
      neg_av_2_26_port, neg_av_2_25_port, neg_av_2_24_port, neg_av_2_23_port, 
      neg_av_2_22_port, neg_av_2_21_port, neg_av_2_20_port, neg_av_2_19_port, 
      neg_av_2_18_port, neg_av_2_17_port, neg_av_2_16_port, neg_av_2_15_port, 
      neg_av_2_14_port, neg_av_2_13_port, neg_av_2_12_port, neg_av_2_11_port, 
      neg_av_2_10_port, neg_av_2_9_port, neg_av_2_8_port, neg_av_2_7_port, 
      neg_av_2_6_port, neg_av_2_5_port, neg_av_2_4_port, neg_av_2_3_port, 
      neg_av_2_2_port, neg_av_2_1_port, neg_av_2_0_port, neg_av_1_31_port, 
      neg_av_1_30_port, neg_av_1_29_port, neg_av_1_28_port, neg_av_1_27_port, 
      neg_av_1_26_port, neg_av_1_25_port, neg_av_1_24_port, neg_av_1_23_port, 
      neg_av_1_22_port, neg_av_1_21_port, neg_av_1_20_port, neg_av_1_19_port, 
      neg_av_1_18_port, neg_av_1_17_port, neg_av_1_16_port, neg_av_1_15_port, 
      neg_av_1_14_port, neg_av_1_13_port, neg_av_1_12_port, neg_av_1_11_port, 
      neg_av_1_10_port, neg_av_1_9_port, neg_av_1_8_port, neg_av_1_7_port, 
      neg_av_1_6_port, neg_av_1_5_port, neg_av_1_4_port, neg_av_1_3_port, 
      neg_av_1_2_port, neg_av_1_1_port, neg_av_1_0_port, neg_av_0_31_port, 
      neg_av_0_30_port, neg_av_0_29_port, neg_av_0_28_port, neg_av_0_27_port, 
      neg_av_0_26_port, neg_av_0_25_port, neg_av_0_24_port, neg_av_0_23_port, 
      neg_av_0_22_port, neg_av_0_21_port, neg_av_0_20_port, neg_av_0_19_port, 
      neg_av_0_18_port, neg_av_0_17_port, neg_av_0_16_port, neg_av_0_15_port, 
      neg_av_0_14_port, neg_av_0_13_port, neg_av_0_12_port, neg_av_0_11_port, 
      neg_av_0_10_port, neg_av_0_9_port, neg_av_0_8_port, neg_av_0_7_port, 
      neg_av_0_6_port, neg_av_0_5_port, neg_av_0_4_port, neg_av_0_3_port, 
      neg_av_0_2_port, neg_av_0_1_port, neg_av_0_0_port, pos_av_7_31_port, 
      pos_av_7_30_port, pos_av_7_29_port, pos_av_7_28_port, pos_av_7_27_port, 
      pos_av_7_26_port, pos_av_7_25_port, pos_av_7_24_port, pos_av_7_23_port, 
      pos_av_7_22_port, pos_av_7_21_port, pos_av_7_20_port, pos_av_7_19_port, 
      pos_av_7_18_port, pos_av_7_17_port, pos_av_7_16_port, pos_av_7_15_port, 
      pos_av_7_14_port, pos_av_7_13_port, pos_av_7_12_port, pos_av_7_11_port, 
      pos_av_7_10_port, pos_av_7_9_port, pos_av_7_8_port, pos_av_7_7_port, 
      pos_av_7_6_port, pos_av_7_5_port, pos_av_7_4_port, pos_av_7_3_port, 
      pos_av_7_2_port, pos_av_7_1_port, pos_av_7_0_port, pos_av_6_31_port, 
      pos_av_6_30_port, pos_av_6_29_port, pos_av_6_28_port, pos_av_6_27_port, 
      pos_av_6_26_port, pos_av_6_25_port, pos_av_6_24_port, pos_av_6_23_port, 
      pos_av_6_22_port, pos_av_6_21_port, pos_av_6_20_port, pos_av_6_19_port, 
      pos_av_6_18_port, pos_av_6_17_port, pos_av_6_16_port, pos_av_6_15_port, 
      pos_av_6_14_port, pos_av_6_13_port, pos_av_6_12_port, pos_av_6_11_port, 
      pos_av_6_10_port, pos_av_6_9_port, pos_av_6_8_port, pos_av_6_7_port, 
      pos_av_6_6_port, pos_av_6_5_port, pos_av_6_4_port, pos_av_6_3_port, 
      pos_av_6_2_port, pos_av_6_1_port, pos_av_6_0_port, pos_av_5_31_port, 
      pos_av_5_30_port, pos_av_5_29_port, pos_av_5_28_port, pos_av_5_27_port, 
      pos_av_5_26_port, pos_av_5_25_port, pos_av_5_24_port, pos_av_5_23_port, 
      pos_av_5_22_port, pos_av_5_21_port, pos_av_5_20_port, pos_av_5_19_port, 
      pos_av_5_18_port, pos_av_5_17_port, pos_av_5_16_port, pos_av_5_15_port, 
      pos_av_5_14_port, pos_av_5_13_port, pos_av_5_12_port, pos_av_5_11_port, 
      pos_av_5_10_port, pos_av_5_9_port, pos_av_5_8_port, pos_av_5_7_port, 
      pos_av_5_6_port, pos_av_5_5_port, pos_av_5_4_port, pos_av_5_3_port, 
      pos_av_5_2_port, pos_av_5_1_port, pos_av_5_0_port, pos_av_4_31_port, 
      pos_av_4_30_port, pos_av_4_29_port, pos_av_4_28_port, pos_av_4_27_port, 
      pos_av_4_26_port, pos_av_4_25_port, pos_av_4_24_port, pos_av_4_23_port, 
      pos_av_4_22_port, pos_av_4_21_port, pos_av_4_20_port, pos_av_4_19_port, 
      pos_av_4_18_port, pos_av_4_17_port, pos_av_4_16_port, pos_av_4_15_port, 
      pos_av_4_14_port, pos_av_4_13_port, pos_av_4_12_port, pos_av_4_11_port, 
      pos_av_4_10_port, pos_av_4_9_port, pos_av_4_8_port, pos_av_4_7_port, 
      pos_av_4_6_port, pos_av_4_5_port, pos_av_4_4_port, pos_av_4_3_port, 
      pos_av_4_2_port, pos_av_4_1_port, pos_av_4_0_port, pos_av_3_31_port, 
      pos_av_3_30_port, pos_av_3_29_port, pos_av_3_28_port, pos_av_3_27_port, 
      pos_av_3_26_port, pos_av_3_25_port, pos_av_3_24_port, pos_av_3_23_port, 
      pos_av_3_22_port, pos_av_3_21_port, pos_av_3_20_port, pos_av_3_19_port, 
      pos_av_3_18_port, pos_av_3_17_port, pos_av_3_16_port, pos_av_3_15_port, 
      pos_av_3_14_port, pos_av_3_13_port, pos_av_3_12_port, pos_av_3_11_port, 
      pos_av_3_10_port, pos_av_3_9_port, pos_av_3_8_port, pos_av_3_7_port, 
      pos_av_3_6_port, pos_av_3_5_port, pos_av_3_4_port, pos_av_3_3_port, 
      pos_av_3_2_port, pos_av_3_1_port, pos_av_3_0_port, pos_av_2_31_port, 
      pos_av_2_30_port, pos_av_2_29_port, pos_av_2_28_port, pos_av_2_27_port, 
      pos_av_2_26_port, pos_av_2_25_port, pos_av_2_24_port, pos_av_2_23_port, 
      pos_av_2_22_port, pos_av_2_21_port, pos_av_2_20_port, pos_av_2_19_port, 
      pos_av_2_18_port, pos_av_2_17_port, pos_av_2_16_port, pos_av_2_15_port, 
      pos_av_2_14_port, pos_av_2_13_port, pos_av_2_12_port, pos_av_2_11_port, 
      pos_av_2_10_port, pos_av_2_9_port, pos_av_2_8_port, pos_av_2_7_port, 
      pos_av_2_6_port, pos_av_2_5_port, pos_av_2_4_port, pos_av_2_3_port, 
      pos_av_2_2_port, pos_av_2_1_port, pos_av_2_0_port, pos_av_1_31_port, 
      pos_av_1_30_port, pos_av_1_29_port, pos_av_1_28_port, pos_av_1_27_port, 
      pos_av_1_26_port, pos_av_1_25_port, pos_av_1_24_port, pos_av_1_23_port, 
      pos_av_1_22_port, pos_av_1_21_port, pos_av_1_20_port, pos_av_1_19_port, 
      pos_av_1_18_port, pos_av_1_17_port, pos_av_1_16_port, pos_av_1_15_port, 
      pos_av_1_14_port, pos_av_1_13_port, pos_av_1_12_port, pos_av_1_11_port, 
      pos_av_1_10_port, pos_av_1_9_port, pos_av_1_8_port, pos_av_1_7_port, 
      pos_av_1_6_port, pos_av_1_5_port, pos_av_1_4_port, pos_av_1_3_port, 
      pos_av_1_2_port, pos_av_1_1_port, pos_av_1_0_port, pos_av_0_31_port, 
      pos_av_0_30_port, pos_av_0_29_port, pos_av_0_28_port, pos_av_0_27_port, 
      pos_av_0_26_port, pos_av_0_25_port, pos_av_0_24_port, pos_av_0_23_port, 
      pos_av_0_22_port, pos_av_0_21_port, pos_av_0_20_port, pos_av_0_19_port, 
      pos_av_0_18_port, pos_av_0_17_port, pos_av_0_16_port, pos_av_0_15_port, 
      pos_av_0_14_port, pos_av_0_13_port, pos_av_0_12_port, pos_av_0_11_port, 
      pos_av_0_10_port, pos_av_0_9_port, pos_av_0_8_port, pos_av_0_7_port, 
      pos_av_0_6_port, pos_av_0_5_port, pos_av_0_4_port, pos_av_0_3_port, 
      pos_av_0_2_port, pos_av_0_1_port, pos_av_0_0_port, sum_vector_13_31_port,
      sum_vector_13_30_port, sum_vector_13_29_port, sum_vector_13_28_port, 
      sum_vector_13_27_port, sum_vector_13_26_port, sum_vector_13_25_port, 
      sum_vector_13_24_port, sum_vector_13_23_port, sum_vector_13_22_port, 
      sum_vector_13_21_port, sum_vector_13_20_port, sum_vector_13_19_port, 
      sum_vector_13_18_port, sum_vector_13_17_port, sum_vector_13_16_port, 
      sum_vector_13_15_port, sum_vector_13_14_port, sum_vector_13_13_port, 
      sum_vector_13_12_port, sum_vector_13_11_port, sum_vector_13_10_port, 
      sum_vector_13_9_port, sum_vector_13_8_port, sum_vector_13_7_port, 
      sum_vector_13_6_port, sum_vector_13_5_port, sum_vector_13_4_port, 
      sum_vector_13_3_port, sum_vector_13_2_port, sum_vector_13_1_port, 
      sum_vector_13_0_port, sum_vector_12_31_port, sum_vector_12_30_port, 
      sum_vector_12_29_port, sum_vector_12_28_port, sum_vector_12_27_port, 
      sum_vector_12_26_port, sum_vector_12_25_port, sum_vector_12_24_port, 
      sum_vector_12_23_port, sum_vector_12_22_port, sum_vector_12_21_port, 
      sum_vector_12_20_port, sum_vector_12_19_port, sum_vector_12_18_port, 
      sum_vector_12_17_port, sum_vector_12_16_port, sum_vector_12_15_port, 
      sum_vector_12_14_port, sum_vector_12_13_port, sum_vector_12_12_port, 
      sum_vector_12_11_port, sum_vector_12_10_port, sum_vector_12_9_port, 
      sum_vector_12_8_port, sum_vector_12_7_port, sum_vector_12_6_port, 
      sum_vector_12_5_port, sum_vector_12_4_port, sum_vector_12_3_port, 
      sum_vector_12_2_port, sum_vector_12_1_port, sum_vector_12_0_port, 
      sum_vector_11_31_port, sum_vector_11_30_port, sum_vector_11_29_port, 
      sum_vector_11_28_port, sum_vector_11_27_port, sum_vector_11_26_port, 
      sum_vector_11_25_port, sum_vector_11_24_port, sum_vector_11_23_port, 
      sum_vector_11_22_port, sum_vector_11_21_port, sum_vector_11_20_port, 
      sum_vector_11_19_port, sum_vector_11_18_port, sum_vector_11_17_port, 
      sum_vector_11_16_port, sum_vector_11_15_port, sum_vector_11_14_port, 
      sum_vector_11_13_port, sum_vector_11_12_port, sum_vector_11_11_port, 
      sum_vector_11_10_port, sum_vector_11_9_port, sum_vector_11_8_port, 
      sum_vector_11_7_port, sum_vector_11_6_port, sum_vector_11_5_port, 
      sum_vector_11_4_port, sum_vector_11_3_port, sum_vector_11_2_port, 
      sum_vector_11_1_port, sum_vector_11_0_port, sum_vector_10_31_port, 
      sum_vector_10_30_port, sum_vector_10_29_port, sum_vector_10_28_port, 
      sum_vector_10_27_port, sum_vector_10_26_port, sum_vector_10_25_port, 
      sum_vector_10_24_port, sum_vector_10_23_port, sum_vector_10_22_port, 
      sum_vector_10_21_port, sum_vector_10_20_port, sum_vector_10_19_port, 
      sum_vector_10_18_port, sum_vector_10_17_port, sum_vector_10_16_port, 
      sum_vector_10_15_port, sum_vector_10_14_port, sum_vector_10_13_port, 
      sum_vector_10_12_port, sum_vector_10_11_port, sum_vector_10_10_port, 
      sum_vector_10_9_port, sum_vector_10_8_port, sum_vector_10_7_port, 
      sum_vector_10_6_port, sum_vector_10_5_port, sum_vector_10_4_port, 
      sum_vector_10_3_port, sum_vector_10_2_port, sum_vector_10_1_port, 
      sum_vector_10_0_port, sum_vector_9_31_port, sum_vector_9_30_port, 
      sum_vector_9_29_port, sum_vector_9_28_port, sum_vector_9_27_port, 
      sum_vector_9_26_port, sum_vector_9_25_port, sum_vector_9_24_port, 
      sum_vector_9_23_port, sum_vector_9_22_port, sum_vector_9_21_port, 
      sum_vector_9_20_port, sum_vector_9_19_port, sum_vector_9_18_port, 
      sum_vector_9_17_port, sum_vector_9_16_port, sum_vector_9_15_port, 
      sum_vector_9_14_port, sum_vector_9_13_port, sum_vector_9_12_port, 
      sum_vector_9_11_port, sum_vector_9_10_port, sum_vector_9_9_port, 
      sum_vector_9_8_port, sum_vector_9_7_port, sum_vector_9_6_port, 
      sum_vector_9_5_port, sum_vector_9_4_port, sum_vector_9_3_port, 
      sum_vector_9_2_port, sum_vector_9_1_port, sum_vector_9_0_port, 
      sum_vector_8_31_port, sum_vector_8_30_port, sum_vector_8_29_port, 
      sum_vector_8_28_port, sum_vector_8_27_port, sum_vector_8_26_port, 
      sum_vector_8_25_port, sum_vector_8_24_port, sum_vector_8_23_port, 
      sum_vector_8_22_port, sum_vector_8_21_port, sum_vector_8_20_port, 
      sum_vector_8_19_port, sum_vector_8_18_port, sum_vector_8_17_port, 
      sum_vector_8_16_port, sum_vector_8_15_port, sum_vector_8_14_port, 
      sum_vector_8_13_port, sum_vector_8_12_port, sum_vector_8_11_port, 
      sum_vector_8_10_port, sum_vector_8_9_port, sum_vector_8_8_port, 
      sum_vector_8_7_port, sum_vector_8_6_port, sum_vector_8_5_port, 
      sum_vector_8_4_port, sum_vector_8_3_port, sum_vector_8_2_port, 
      sum_vector_8_1_port, sum_vector_8_0_port, sum_vector_7_31_port, 
      sum_vector_7_30_port, sum_vector_7_29_port, sum_vector_7_28_port, 
      sum_vector_7_27_port, sum_vector_7_26_port, sum_vector_7_25_port, 
      sum_vector_7_24_port, sum_vector_7_23_port, sum_vector_7_22_port, 
      sum_vector_7_21_port, sum_vector_7_20_port, sum_vector_7_19_port, 
      sum_vector_7_18_port, sum_vector_7_17_port, sum_vector_7_16_port, 
      sum_vector_7_15_port, sum_vector_7_14_port, sum_vector_7_13_port, 
      sum_vector_7_12_port, sum_vector_7_11_port, sum_vector_7_10_port, 
      sum_vector_7_9_port, sum_vector_7_8_port, sum_vector_7_7_port, 
      sum_vector_7_6_port, sum_vector_7_5_port, sum_vector_7_4_port, 
      sum_vector_7_3_port, sum_vector_7_2_port, sum_vector_7_1_port, 
      sum_vector_7_0_port, sum_vector_6_31_port, sum_vector_6_30_port, 
      sum_vector_6_29_port, sum_vector_6_28_port, sum_vector_6_27_port, 
      sum_vector_6_26_port, sum_vector_6_25_port, sum_vector_6_24_port, 
      sum_vector_6_23_port, sum_vector_6_22_port, sum_vector_6_21_port, 
      sum_vector_6_20_port, sum_vector_6_19_port, sum_vector_6_18_port, 
      sum_vector_6_17_port, sum_vector_6_16_port, sum_vector_6_15_port, 
      sum_vector_6_14_port, sum_vector_6_13_port, sum_vector_6_12_port, 
      sum_vector_6_11_port, sum_vector_6_10_port, sum_vector_6_9_port, 
      sum_vector_6_8_port, sum_vector_6_7_port, sum_vector_6_6_port, 
      sum_vector_6_5_port, sum_vector_6_4_port, sum_vector_6_3_port, 
      sum_vector_6_2_port, sum_vector_6_1_port, sum_vector_6_0_port, 
      sum_vector_5_31_port, sum_vector_5_30_port, sum_vector_5_29_port, 
      sum_vector_5_28_port, sum_vector_5_27_port, sum_vector_5_26_port, 
      sum_vector_5_25_port, sum_vector_5_24_port, sum_vector_5_23_port, 
      sum_vector_5_22_port, sum_vector_5_21_port, sum_vector_5_20_port, 
      sum_vector_5_19_port, sum_vector_5_18_port, sum_vector_5_17_port, 
      sum_vector_5_16_port, sum_vector_5_15_port, sum_vector_5_14_port, 
      sum_vector_5_13_port, sum_vector_5_12_port, sum_vector_5_11_port, 
      sum_vector_5_10_port, sum_vector_5_9_port, sum_vector_5_8_port, 
      sum_vector_5_7_port, sum_vector_5_6_port, sum_vector_5_5_port, 
      sum_vector_5_4_port, sum_vector_5_3_port, sum_vector_5_2_port, 
      sum_vector_5_1_port, sum_vector_5_0_port, sum_vector_4_31_port, 
      sum_vector_4_30_port, sum_vector_4_29_port, sum_vector_4_28_port, 
      sum_vector_4_27_port, sum_vector_4_26_port, sum_vector_4_25_port, 
      sum_vector_4_24_port, sum_vector_4_23_port, sum_vector_4_22_port, 
      sum_vector_4_21_port, sum_vector_4_20_port, sum_vector_4_19_port, 
      sum_vector_4_18_port, sum_vector_4_17_port, sum_vector_4_16_port, 
      sum_vector_4_15_port, sum_vector_4_14_port, sum_vector_4_13_port, 
      sum_vector_4_12_port, sum_vector_4_11_port, sum_vector_4_10_port, 
      sum_vector_4_9_port, sum_vector_4_8_port, sum_vector_4_7_port, 
      sum_vector_4_6_port, sum_vector_4_5_port, sum_vector_4_4_port, 
      sum_vector_4_3_port, sum_vector_4_2_port, sum_vector_4_1_port, 
      sum_vector_4_0_port, sum_vector_3_31_port, sum_vector_3_30_port, 
      sum_vector_3_29_port, sum_vector_3_28_port, sum_vector_3_27_port, 
      sum_vector_3_26_port, sum_vector_3_25_port, sum_vector_3_24_port, 
      sum_vector_3_23_port, sum_vector_3_22_port, sum_vector_3_21_port, 
      sum_vector_3_20_port, sum_vector_3_19_port, sum_vector_3_18_port, 
      sum_vector_3_17_port, sum_vector_3_16_port, sum_vector_3_15_port, 
      sum_vector_3_14_port, sum_vector_3_13_port, sum_vector_3_12_port, 
      sum_vector_3_11_port, sum_vector_3_10_port, sum_vector_3_9_port, 
      sum_vector_3_8_port, sum_vector_3_7_port, sum_vector_3_6_port, 
      sum_vector_3_5_port, sum_vector_3_4_port, sum_vector_3_3_port, 
      sum_vector_3_2_port, sum_vector_3_1_port, sum_vector_3_0_port, 
      sum_vector_2_31_port, sum_vector_2_30_port, sum_vector_2_29_port, 
      sum_vector_2_28_port, sum_vector_2_27_port, sum_vector_2_26_port, 
      sum_vector_2_25_port, sum_vector_2_24_port, sum_vector_2_23_port, 
      sum_vector_2_22_port, sum_vector_2_21_port, sum_vector_2_20_port, 
      sum_vector_2_19_port, sum_vector_2_18_port, sum_vector_2_17_port, 
      sum_vector_2_16_port, sum_vector_2_15_port, sum_vector_2_14_port, 
      sum_vector_2_13_port, sum_vector_2_12_port, sum_vector_2_11_port, 
      sum_vector_2_10_port, sum_vector_2_9_port, sum_vector_2_8_port, 
      sum_vector_2_7_port, sum_vector_2_6_port, sum_vector_2_5_port, 
      sum_vector_2_4_port, sum_vector_2_3_port, sum_vector_2_2_port, 
      sum_vector_2_1_port, sum_vector_2_0_port, sum_vector_1_31_port, 
      sum_vector_1_30_port, sum_vector_1_29_port, sum_vector_1_28_port, 
      sum_vector_1_27_port, sum_vector_1_26_port, sum_vector_1_25_port, 
      sum_vector_1_24_port, sum_vector_1_23_port, sum_vector_1_22_port, 
      sum_vector_1_21_port, sum_vector_1_20_port, sum_vector_1_19_port, 
      sum_vector_1_18_port, sum_vector_1_17_port, sum_vector_1_16_port, 
      sum_vector_1_15_port, sum_vector_1_14_port, sum_vector_1_13_port, 
      sum_vector_1_12_port, sum_vector_1_11_port, sum_vector_1_10_port, 
      sum_vector_1_9_port, sum_vector_1_8_port, sum_vector_1_7_port, 
      sum_vector_1_6_port, sum_vector_1_5_port, sum_vector_1_4_port, 
      sum_vector_1_3_port, sum_vector_1_2_port, sum_vector_1_1_port, 
      sum_vector_1_0_port, sum_vector_0_31_port, sum_vector_0_30_port, 
      sum_vector_0_29_port, sum_vector_0_28_port, sum_vector_0_27_port, 
      sum_vector_0_26_port, sum_vector_0_25_port, sum_vector_0_24_port, 
      sum_vector_0_23_port, sum_vector_0_22_port, sum_vector_0_21_port, 
      sum_vector_0_20_port, sum_vector_0_19_port, sum_vector_0_18_port, 
      sum_vector_0_17_port, sum_vector_0_16_port, sum_vector_0_15_port, 
      sum_vector_0_14_port, sum_vector_0_13_port, sum_vector_0_12_port, 
      sum_vector_0_11_port, sum_vector_0_10_port, sum_vector_0_9_port, 
      sum_vector_0_8_port, sum_vector_0_7_port, sum_vector_0_6_port, 
      sum_vector_0_5_port, sum_vector_0_4_port, sum_vector_0_3_port, 
      sum_vector_0_2_port, sum_vector_0_1_port, sum_vector_0_0_port, n_1164, 
      n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, 
      n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, 
      n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, 
      n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, 
      n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, 
      n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, 
      n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, 
      n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, 
      n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, 
      n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, 
      n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, 
      n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, 
      n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, 
      n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, 
      n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, 
      n_1408, n_1409, n_1410 : std_logic;

begin
   
   X_Logic0_port <= '0';
   sh0_0 : shift_NBIT32_SHIFT0 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_0_31_port, pos_a(30) => 
                           pos_av_0_30_port, pos_a(29) => pos_av_0_29_port, 
                           pos_a(28) => pos_av_0_28_port, pos_a(27) => 
                           pos_av_0_27_port, pos_a(26) => pos_av_0_26_port, 
                           pos_a(25) => pos_av_0_25_port, pos_a(24) => 
                           pos_av_0_24_port, pos_a(23) => pos_av_0_23_port, 
                           pos_a(22) => pos_av_0_22_port, pos_a(21) => 
                           pos_av_0_21_port, pos_a(20) => pos_av_0_20_port, 
                           pos_a(19) => pos_av_0_19_port, pos_a(18) => 
                           pos_av_0_18_port, pos_a(17) => pos_av_0_17_port, 
                           pos_a(16) => pos_av_0_16_port, pos_a(15) => 
                           pos_av_0_15_port, pos_a(14) => pos_av_0_14_port, 
                           pos_a(13) => pos_av_0_13_port, pos_a(12) => 
                           pos_av_0_12_port, pos_a(11) => pos_av_0_11_port, 
                           pos_a(10) => pos_av_0_10_port, pos_a(9) => 
                           pos_av_0_9_port, pos_a(8) => pos_av_0_8_port, 
                           pos_a(7) => pos_av_0_7_port, pos_a(6) => 
                           pos_av_0_6_port, pos_a(5) => pos_av_0_5_port, 
                           pos_a(4) => pos_av_0_4_port, pos_a(3) => 
                           pos_av_0_3_port, pos_a(2) => pos_av_0_2_port, 
                           pos_a(1) => pos_av_0_1_port, pos_a(0) => 
                           pos_av_0_0_port, neg_a(31) => neg_av_0_31_port, 
                           neg_a(30) => neg_av_0_30_port, neg_a(29) => 
                           neg_av_0_29_port, neg_a(28) => neg_av_0_28_port, 
                           neg_a(27) => neg_av_0_27_port, neg_a(26) => 
                           neg_av_0_26_port, neg_a(25) => neg_av_0_25_port, 
                           neg_a(24) => neg_av_0_24_port, neg_a(23) => 
                           neg_av_0_23_port, neg_a(22) => neg_av_0_22_port, 
                           neg_a(21) => neg_av_0_21_port, neg_a(20) => 
                           neg_av_0_20_port, neg_a(19) => neg_av_0_19_port, 
                           neg_a(18) => neg_av_0_18_port, neg_a(17) => 
                           neg_av_0_17_port, neg_a(16) => neg_av_0_16_port, 
                           neg_a(15) => neg_av_0_15_port, neg_a(14) => 
                           neg_av_0_14_port, neg_a(13) => neg_av_0_13_port, 
                           neg_a(12) => neg_av_0_12_port, neg_a(11) => 
                           neg_av_0_11_port, neg_a(10) => neg_av_0_10_port, 
                           neg_a(9) => neg_av_0_9_port, neg_a(8) => 
                           neg_av_0_8_port, neg_a(7) => neg_av_0_7_port, 
                           neg_a(6) => neg_av_0_6_port, neg_a(5) => 
                           neg_av_0_5_port, neg_a(4) => neg_av_0_4_port, 
                           neg_a(3) => neg_av_0_3_port, neg_a(2) => 
                           neg_av_0_2_port, neg_a(1) => neg_av_0_1_port, 
                           neg_a(0) => neg_av_0_0_port, pos_2a(31) => 
                           pos_2av_0_31_port, pos_2a(30) => pos_2av_0_30_port, 
                           pos_2a(29) => pos_2av_0_29_port, pos_2a(28) => 
                           pos_2av_0_28_port, pos_2a(27) => pos_2av_0_27_port, 
                           pos_2a(26) => pos_2av_0_26_port, pos_2a(25) => 
                           pos_2av_0_25_port, pos_2a(24) => pos_2av_0_24_port, 
                           pos_2a(23) => pos_2av_0_23_port, pos_2a(22) => 
                           pos_2av_0_22_port, pos_2a(21) => pos_2av_0_21_port, 
                           pos_2a(20) => pos_2av_0_20_port, pos_2a(19) => 
                           pos_2av_0_19_port, pos_2a(18) => pos_2av_0_18_port, 
                           pos_2a(17) => pos_2av_0_17_port, pos_2a(16) => 
                           pos_2av_0_16_port, pos_2a(15) => pos_2av_0_15_port, 
                           pos_2a(14) => pos_2av_0_14_port, pos_2a(13) => 
                           pos_2av_0_13_port, pos_2a(12) => pos_2av_0_12_port, 
                           pos_2a(11) => pos_2av_0_11_port, pos_2a(10) => 
                           pos_2av_0_10_port, pos_2a(9) => pos_2av_0_9_port, 
                           pos_2a(8) => pos_2av_0_8_port, pos_2a(7) => 
                           pos_2av_0_7_port, pos_2a(6) => pos_2av_0_6_port, 
                           pos_2a(5) => pos_2av_0_5_port, pos_2a(4) => 
                           pos_2av_0_4_port, pos_2a(3) => pos_2av_0_3_port, 
                           pos_2a(2) => pos_2av_0_2_port, pos_2a(1) => 
                           pos_2av_0_1_port, pos_2a(0) => n_1164, neg_2a(31) =>
                           neg_2av_0_31_port, neg_2a(30) => neg_2av_0_30_port, 
                           neg_2a(29) => neg_2av_0_29_port, neg_2a(28) => 
                           neg_2av_0_28_port, neg_2a(27) => neg_2av_0_27_port, 
                           neg_2a(26) => neg_2av_0_26_port, neg_2a(25) => 
                           neg_2av_0_25_port, neg_2a(24) => neg_2av_0_24_port, 
                           neg_2a(23) => neg_2av_0_23_port, neg_2a(22) => 
                           neg_2av_0_22_port, neg_2a(21) => neg_2av_0_21_port, 
                           neg_2a(20) => neg_2av_0_20_port, neg_2a(19) => 
                           neg_2av_0_19_port, neg_2a(18) => neg_2av_0_18_port, 
                           neg_2a(17) => neg_2av_0_17_port, neg_2a(16) => 
                           neg_2av_0_16_port, neg_2a(15) => neg_2av_0_15_port, 
                           neg_2a(14) => neg_2av_0_14_port, neg_2a(13) => 
                           neg_2av_0_13_port, neg_2a(12) => neg_2av_0_12_port, 
                           neg_2a(11) => neg_2av_0_11_port, neg_2a(10) => 
                           neg_2av_0_10_port, neg_2a(9) => neg_2av_0_9_port, 
                           neg_2a(8) => neg_2av_0_8_port, neg_2a(7) => 
                           neg_2av_0_7_port, neg_2a(6) => neg_2av_0_6_port, 
                           neg_2a(5) => neg_2av_0_5_port, neg_2a(4) => 
                           neg_2av_0_4_port, neg_2a(3) => neg_2av_0_3_port, 
                           neg_2a(2) => neg_2av_0_2_port, neg_2a(1) => 
                           neg_2av_0_1_port, neg_2a(0) => n_1165);
   vp0_0 : vp_NBIT32_0 port map( pos_a(31) => pos_av_0_31_port, pos_a(30) => 
                           pos_av_0_30_port, pos_a(29) => pos_av_0_29_port, 
                           pos_a(28) => pos_av_0_28_port, pos_a(27) => 
                           pos_av_0_27_port, pos_a(26) => pos_av_0_26_port, 
                           pos_a(25) => pos_av_0_25_port, pos_a(24) => 
                           pos_av_0_24_port, pos_a(23) => pos_av_0_23_port, 
                           pos_a(22) => pos_av_0_22_port, pos_a(21) => 
                           pos_av_0_21_port, pos_a(20) => pos_av_0_20_port, 
                           pos_a(19) => pos_av_0_19_port, pos_a(18) => 
                           pos_av_0_18_port, pos_a(17) => pos_av_0_17_port, 
                           pos_a(16) => pos_av_0_16_port, pos_a(15) => 
                           pos_av_0_15_port, pos_a(14) => pos_av_0_14_port, 
                           pos_a(13) => pos_av_0_13_port, pos_a(12) => 
                           pos_av_0_12_port, pos_a(11) => pos_av_0_11_port, 
                           pos_a(10) => pos_av_0_10_port, pos_a(9) => 
                           pos_av_0_9_port, pos_a(8) => pos_av_0_8_port, 
                           pos_a(7) => pos_av_0_7_port, pos_a(6) => 
                           pos_av_0_6_port, pos_a(5) => pos_av_0_5_port, 
                           pos_a(4) => pos_av_0_4_port, pos_a(3) => 
                           pos_av_0_3_port, pos_a(2) => pos_av_0_2_port, 
                           pos_a(1) => pos_av_0_1_port, pos_a(0) => 
                           pos_av_0_0_port, neg_a(31) => neg_av_0_31_port, 
                           neg_a(30) => neg_av_0_30_port, neg_a(29) => 
                           neg_av_0_29_port, neg_a(28) => neg_av_0_28_port, 
                           neg_a(27) => neg_av_0_27_port, neg_a(26) => 
                           neg_av_0_26_port, neg_a(25) => neg_av_0_25_port, 
                           neg_a(24) => neg_av_0_24_port, neg_a(23) => 
                           neg_av_0_23_port, neg_a(22) => neg_av_0_22_port, 
                           neg_a(21) => neg_av_0_21_port, neg_a(20) => 
                           neg_av_0_20_port, neg_a(19) => neg_av_0_19_port, 
                           neg_a(18) => neg_av_0_18_port, neg_a(17) => 
                           neg_av_0_17_port, neg_a(16) => neg_av_0_16_port, 
                           neg_a(15) => neg_av_0_15_port, neg_a(14) => 
                           neg_av_0_14_port, neg_a(13) => neg_av_0_13_port, 
                           neg_a(12) => neg_av_0_12_port, neg_a(11) => 
                           neg_av_0_11_port, neg_a(10) => neg_av_0_10_port, 
                           neg_a(9) => neg_av_0_9_port, neg_a(8) => 
                           neg_av_0_8_port, neg_a(7) => neg_av_0_7_port, 
                           neg_a(6) => neg_av_0_6_port, neg_a(5) => 
                           neg_av_0_5_port, neg_a(4) => neg_av_0_4_port, 
                           neg_a(3) => neg_av_0_3_port, neg_a(2) => 
                           neg_av_0_2_port, neg_a(1) => neg_av_0_1_port, 
                           neg_a(0) => neg_av_0_0_port, pos_2a(31) => 
                           pos_2av_0_31_port, pos_2a(30) => pos_2av_0_30_port, 
                           pos_2a(29) => pos_2av_0_29_port, pos_2a(28) => 
                           pos_2av_0_28_port, pos_2a(27) => pos_2av_0_27_port, 
                           pos_2a(26) => pos_2av_0_26_port, pos_2a(25) => 
                           pos_2av_0_25_port, pos_2a(24) => pos_2av_0_24_port, 
                           pos_2a(23) => pos_2av_0_23_port, pos_2a(22) => 
                           pos_2av_0_22_port, pos_2a(21) => pos_2av_0_21_port, 
                           pos_2a(20) => pos_2av_0_20_port, pos_2a(19) => 
                           pos_2av_0_19_port, pos_2a(18) => pos_2av_0_18_port, 
                           pos_2a(17) => pos_2av_0_17_port, pos_2a(16) => 
                           pos_2av_0_16_port, pos_2a(15) => pos_2av_0_15_port, 
                           pos_2a(14) => pos_2av_0_14_port, pos_2a(13) => 
                           pos_2av_0_13_port, pos_2a(12) => pos_2av_0_12_port, 
                           pos_2a(11) => pos_2av_0_11_port, pos_2a(10) => 
                           pos_2av_0_10_port, pos_2a(9) => pos_2av_0_9_port, 
                           pos_2a(8) => pos_2av_0_8_port, pos_2a(7) => 
                           pos_2av_0_7_port, pos_2a(6) => pos_2av_0_6_port, 
                           pos_2a(5) => pos_2av_0_5_port, pos_2a(4) => 
                           pos_2av_0_4_port, pos_2a(3) => pos_2av_0_3_port, 
                           pos_2a(2) => pos_2av_0_2_port, pos_2a(1) => 
                           pos_2av_0_1_port, pos_2a(0) => pos_2av_0_0_port, 
                           neg_2a(31) => neg_2av_0_31_port, neg_2a(30) => 
                           neg_2av_0_30_port, neg_2a(29) => neg_2av_0_29_port, 
                           neg_2a(28) => neg_2av_0_28_port, neg_2a(27) => 
                           neg_2av_0_27_port, neg_2a(26) => neg_2av_0_26_port, 
                           neg_2a(25) => neg_2av_0_25_port, neg_2a(24) => 
                           neg_2av_0_24_port, neg_2a(23) => neg_2av_0_23_port, 
                           neg_2a(22) => neg_2av_0_22_port, neg_2a(21) => 
                           neg_2av_0_21_port, neg_2a(20) => neg_2av_0_20_port, 
                           neg_2a(19) => neg_2av_0_19_port, neg_2a(18) => 
                           neg_2av_0_18_port, neg_2a(17) => neg_2av_0_17_port, 
                           neg_2a(16) => neg_2av_0_16_port, neg_2a(15) => 
                           neg_2av_0_15_port, neg_2a(14) => neg_2av_0_14_port, 
                           neg_2a(13) => neg_2av_0_13_port, neg_2a(12) => 
                           neg_2av_0_12_port, neg_2a(11) => neg_2av_0_11_port, 
                           neg_2a(10) => neg_2av_0_10_port, neg_2a(9) => 
                           neg_2av_0_9_port, neg_2a(8) => neg_2av_0_8_port, 
                           neg_2a(7) => neg_2av_0_7_port, neg_2a(6) => 
                           neg_2av_0_6_port, neg_2a(5) => neg_2av_0_5_port, 
                           neg_2a(4) => neg_2av_0_4_port, neg_2a(3) => 
                           neg_2av_0_3_port, neg_2a(2) => neg_2av_0_2_port, 
                           neg_2a(1) => neg_2av_0_1_port, neg_2a(0) => 
                           neg_2av_0_0_port, sel(2) => b(1), sel(1) => b(0), 
                           sel(0) => X_Logic0_port, s_out(31) => 
                           sum_vector_0_31_port, s_out(30) => 
                           sum_vector_0_30_port, s_out(29) => 
                           sum_vector_0_29_port, s_out(28) => 
                           sum_vector_0_28_port, s_out(27) => 
                           sum_vector_0_27_port, s_out(26) => 
                           sum_vector_0_26_port, s_out(25) => 
                           sum_vector_0_25_port, s_out(24) => 
                           sum_vector_0_24_port, s_out(23) => 
                           sum_vector_0_23_port, s_out(22) => 
                           sum_vector_0_22_port, s_out(21) => 
                           sum_vector_0_21_port, s_out(20) => 
                           sum_vector_0_20_port, s_out(19) => 
                           sum_vector_0_19_port, s_out(18) => 
                           sum_vector_0_18_port, s_out(17) => 
                           sum_vector_0_17_port, s_out(16) => 
                           sum_vector_0_16_port, s_out(15) => 
                           sum_vector_0_15_port, s_out(14) => 
                           sum_vector_0_14_port, s_out(13) => 
                           sum_vector_0_13_port, s_out(12) => 
                           sum_vector_0_12_port, s_out(11) => 
                           sum_vector_0_11_port, s_out(10) => 
                           sum_vector_0_10_port, s_out(9) => 
                           sum_vector_0_9_port, s_out(8) => sum_vector_0_8_port
                           , s_out(7) => sum_vector_0_7_port, s_out(6) => 
                           sum_vector_0_6_port, s_out(5) => sum_vector_0_5_port
                           , s_out(4) => sum_vector_0_4_port, s_out(3) => 
                           sum_vector_0_3_port, s_out(2) => sum_vector_0_2_port
                           , s_out(1) => sum_vector_0_1_port, s_out(0) => 
                           sum_vector_0_0_port);
   sh1_1 : shift_NBIT32_SHIFT1 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_1_31_port, pos_a(30) => 
                           pos_av_1_30_port, pos_a(29) => pos_av_1_29_port, 
                           pos_a(28) => pos_av_1_28_port, pos_a(27) => 
                           pos_av_1_27_port, pos_a(26) => pos_av_1_26_port, 
                           pos_a(25) => pos_av_1_25_port, pos_a(24) => 
                           pos_av_1_24_port, pos_a(23) => pos_av_1_23_port, 
                           pos_a(22) => pos_av_1_22_port, pos_a(21) => 
                           pos_av_1_21_port, pos_a(20) => pos_av_1_20_port, 
                           pos_a(19) => pos_av_1_19_port, pos_a(18) => 
                           pos_av_1_18_port, pos_a(17) => pos_av_1_17_port, 
                           pos_a(16) => pos_av_1_16_port, pos_a(15) => 
                           pos_av_1_15_port, pos_a(14) => pos_av_1_14_port, 
                           pos_a(13) => pos_av_1_13_port, pos_a(12) => 
                           pos_av_1_12_port, pos_a(11) => pos_av_1_11_port, 
                           pos_a(10) => pos_av_1_10_port, pos_a(9) => 
                           pos_av_1_9_port, pos_a(8) => pos_av_1_8_port, 
                           pos_a(7) => pos_av_1_7_port, pos_a(6) => 
                           pos_av_1_6_port, pos_a(5) => pos_av_1_5_port, 
                           pos_a(4) => pos_av_1_4_port, pos_a(3) => 
                           pos_av_1_3_port, pos_a(2) => pos_av_1_2_port, 
                           pos_a(1) => n_1166, pos_a(0) => n_1167, neg_a(31) =>
                           neg_av_1_31_port, neg_a(30) => neg_av_1_30_port, 
                           neg_a(29) => neg_av_1_29_port, neg_a(28) => 
                           neg_av_1_28_port, neg_a(27) => neg_av_1_27_port, 
                           neg_a(26) => neg_av_1_26_port, neg_a(25) => 
                           neg_av_1_25_port, neg_a(24) => neg_av_1_24_port, 
                           neg_a(23) => neg_av_1_23_port, neg_a(22) => 
                           neg_av_1_22_port, neg_a(21) => neg_av_1_21_port, 
                           neg_a(20) => neg_av_1_20_port, neg_a(19) => 
                           neg_av_1_19_port, neg_a(18) => neg_av_1_18_port, 
                           neg_a(17) => neg_av_1_17_port, neg_a(16) => 
                           neg_av_1_16_port, neg_a(15) => neg_av_1_15_port, 
                           neg_a(14) => neg_av_1_14_port, neg_a(13) => 
                           neg_av_1_13_port, neg_a(12) => neg_av_1_12_port, 
                           neg_a(11) => neg_av_1_11_port, neg_a(10) => 
                           neg_av_1_10_port, neg_a(9) => neg_av_1_9_port, 
                           neg_a(8) => neg_av_1_8_port, neg_a(7) => 
                           neg_av_1_7_port, neg_a(6) => neg_av_1_6_port, 
                           neg_a(5) => neg_av_1_5_port, neg_a(4) => 
                           neg_av_1_4_port, neg_a(3) => neg_av_1_3_port, 
                           neg_a(2) => neg_av_1_2_port, neg_a(1) => n_1168, 
                           neg_a(0) => n_1169, pos_2a(31) => pos_2av_1_31_port,
                           pos_2a(30) => pos_2av_1_30_port, pos_2a(29) => 
                           pos_2av_1_29_port, pos_2a(28) => pos_2av_1_28_port, 
                           pos_2a(27) => pos_2av_1_27_port, pos_2a(26) => 
                           pos_2av_1_26_port, pos_2a(25) => pos_2av_1_25_port, 
                           pos_2a(24) => pos_2av_1_24_port, pos_2a(23) => 
                           pos_2av_1_23_port, pos_2a(22) => pos_2av_1_22_port, 
                           pos_2a(21) => pos_2av_1_21_port, pos_2a(20) => 
                           pos_2av_1_20_port, pos_2a(19) => pos_2av_1_19_port, 
                           pos_2a(18) => pos_2av_1_18_port, pos_2a(17) => 
                           pos_2av_1_17_port, pos_2a(16) => pos_2av_1_16_port, 
                           pos_2a(15) => pos_2av_1_15_port, pos_2a(14) => 
                           pos_2av_1_14_port, pos_2a(13) => pos_2av_1_13_port, 
                           pos_2a(12) => pos_2av_1_12_port, pos_2a(11) => 
                           pos_2av_1_11_port, pos_2a(10) => pos_2av_1_10_port, 
                           pos_2a(9) => pos_2av_1_9_port, pos_2a(8) => 
                           pos_2av_1_8_port, pos_2a(7) => pos_2av_1_7_port, 
                           pos_2a(6) => pos_2av_1_6_port, pos_2a(5) => 
                           pos_2av_1_5_port, pos_2a(4) => pos_2av_1_4_port, 
                           pos_2a(3) => pos_2av_1_3_port, pos_2a(2) => n_1170, 
                           pos_2a(1) => n_1171, pos_2a(0) => n_1172, neg_2a(31)
                           => neg_2av_1_31_port, neg_2a(30) => 
                           neg_2av_1_30_port, neg_2a(29) => neg_2av_1_29_port, 
                           neg_2a(28) => neg_2av_1_28_port, neg_2a(27) => 
                           neg_2av_1_27_port, neg_2a(26) => neg_2av_1_26_port, 
                           neg_2a(25) => neg_2av_1_25_port, neg_2a(24) => 
                           neg_2av_1_24_port, neg_2a(23) => neg_2av_1_23_port, 
                           neg_2a(22) => neg_2av_1_22_port, neg_2a(21) => 
                           neg_2av_1_21_port, neg_2a(20) => neg_2av_1_20_port, 
                           neg_2a(19) => neg_2av_1_19_port, neg_2a(18) => 
                           neg_2av_1_18_port, neg_2a(17) => neg_2av_1_17_port, 
                           neg_2a(16) => neg_2av_1_16_port, neg_2a(15) => 
                           neg_2av_1_15_port, neg_2a(14) => neg_2av_1_14_port, 
                           neg_2a(13) => neg_2av_1_13_port, neg_2a(12) => 
                           neg_2av_1_12_port, neg_2a(11) => neg_2av_1_11_port, 
                           neg_2a(10) => neg_2av_1_10_port, neg_2a(9) => 
                           neg_2av_1_9_port, neg_2a(8) => neg_2av_1_8_port, 
                           neg_2a(7) => neg_2av_1_7_port, neg_2a(6) => 
                           neg_2av_1_6_port, neg_2a(5) => neg_2av_1_5_port, 
                           neg_2a(4) => neg_2av_1_4_port, neg_2a(3) => 
                           neg_2av_1_3_port, neg_2a(2) => n_1173, neg_2a(1) => 
                           n_1174, neg_2a(0) => n_1175);
   vp1_1 : vp_NBIT32_7 port map( pos_a(31) => pos_av_1_31_port, pos_a(30) => 
                           pos_av_1_30_port, pos_a(29) => pos_av_1_29_port, 
                           pos_a(28) => pos_av_1_28_port, pos_a(27) => 
                           pos_av_1_27_port, pos_a(26) => pos_av_1_26_port, 
                           pos_a(25) => pos_av_1_25_port, pos_a(24) => 
                           pos_av_1_24_port, pos_a(23) => pos_av_1_23_port, 
                           pos_a(22) => pos_av_1_22_port, pos_a(21) => 
                           pos_av_1_21_port, pos_a(20) => pos_av_1_20_port, 
                           pos_a(19) => pos_av_1_19_port, pos_a(18) => 
                           pos_av_1_18_port, pos_a(17) => pos_av_1_17_port, 
                           pos_a(16) => pos_av_1_16_port, pos_a(15) => 
                           pos_av_1_15_port, pos_a(14) => pos_av_1_14_port, 
                           pos_a(13) => pos_av_1_13_port, pos_a(12) => 
                           pos_av_1_12_port, pos_a(11) => pos_av_1_11_port, 
                           pos_a(10) => pos_av_1_10_port, pos_a(9) => 
                           pos_av_1_9_port, pos_a(8) => pos_av_1_8_port, 
                           pos_a(7) => pos_av_1_7_port, pos_a(6) => 
                           pos_av_1_6_port, pos_a(5) => pos_av_1_5_port, 
                           pos_a(4) => pos_av_1_4_port, pos_a(3) => 
                           pos_av_1_3_port, pos_a(2) => pos_av_1_2_port, 
                           pos_a(1) => pos_av_1_1_port, pos_a(0) => 
                           pos_av_1_0_port, neg_a(31) => neg_av_1_31_port, 
                           neg_a(30) => neg_av_1_30_port, neg_a(29) => 
                           neg_av_1_29_port, neg_a(28) => neg_av_1_28_port, 
                           neg_a(27) => neg_av_1_27_port, neg_a(26) => 
                           neg_av_1_26_port, neg_a(25) => neg_av_1_25_port, 
                           neg_a(24) => neg_av_1_24_port, neg_a(23) => 
                           neg_av_1_23_port, neg_a(22) => neg_av_1_22_port, 
                           neg_a(21) => neg_av_1_21_port, neg_a(20) => 
                           neg_av_1_20_port, neg_a(19) => neg_av_1_19_port, 
                           neg_a(18) => neg_av_1_18_port, neg_a(17) => 
                           neg_av_1_17_port, neg_a(16) => neg_av_1_16_port, 
                           neg_a(15) => neg_av_1_15_port, neg_a(14) => 
                           neg_av_1_14_port, neg_a(13) => neg_av_1_13_port, 
                           neg_a(12) => neg_av_1_12_port, neg_a(11) => 
                           neg_av_1_11_port, neg_a(10) => neg_av_1_10_port, 
                           neg_a(9) => neg_av_1_9_port, neg_a(8) => 
                           neg_av_1_8_port, neg_a(7) => neg_av_1_7_port, 
                           neg_a(6) => neg_av_1_6_port, neg_a(5) => 
                           neg_av_1_5_port, neg_a(4) => neg_av_1_4_port, 
                           neg_a(3) => neg_av_1_3_port, neg_a(2) => 
                           neg_av_1_2_port, neg_a(1) => neg_av_1_1_port, 
                           neg_a(0) => neg_av_1_0_port, pos_2a(31) => 
                           pos_2av_1_31_port, pos_2a(30) => pos_2av_1_30_port, 
                           pos_2a(29) => pos_2av_1_29_port, pos_2a(28) => 
                           pos_2av_1_28_port, pos_2a(27) => pos_2av_1_27_port, 
                           pos_2a(26) => pos_2av_1_26_port, pos_2a(25) => 
                           pos_2av_1_25_port, pos_2a(24) => pos_2av_1_24_port, 
                           pos_2a(23) => pos_2av_1_23_port, pos_2a(22) => 
                           pos_2av_1_22_port, pos_2a(21) => pos_2av_1_21_port, 
                           pos_2a(20) => pos_2av_1_20_port, pos_2a(19) => 
                           pos_2av_1_19_port, pos_2a(18) => pos_2av_1_18_port, 
                           pos_2a(17) => pos_2av_1_17_port, pos_2a(16) => 
                           pos_2av_1_16_port, pos_2a(15) => pos_2av_1_15_port, 
                           pos_2a(14) => pos_2av_1_14_port, pos_2a(13) => 
                           pos_2av_1_13_port, pos_2a(12) => pos_2av_1_12_port, 
                           pos_2a(11) => pos_2av_1_11_port, pos_2a(10) => 
                           pos_2av_1_10_port, pos_2a(9) => pos_2av_1_9_port, 
                           pos_2a(8) => pos_2av_1_8_port, pos_2a(7) => 
                           pos_2av_1_7_port, pos_2a(6) => pos_2av_1_6_port, 
                           pos_2a(5) => pos_2av_1_5_port, pos_2a(4) => 
                           pos_2av_1_4_port, pos_2a(3) => pos_2av_1_3_port, 
                           pos_2a(2) => pos_2av_1_2_port, pos_2a(1) => 
                           pos_2av_1_1_port, pos_2a(0) => pos_2av_1_0_port, 
                           neg_2a(31) => neg_2av_1_31_port, neg_2a(30) => 
                           neg_2av_1_30_port, neg_2a(29) => neg_2av_1_29_port, 
                           neg_2a(28) => neg_2av_1_28_port, neg_2a(27) => 
                           neg_2av_1_27_port, neg_2a(26) => neg_2av_1_26_port, 
                           neg_2a(25) => neg_2av_1_25_port, neg_2a(24) => 
                           neg_2av_1_24_port, neg_2a(23) => neg_2av_1_23_port, 
                           neg_2a(22) => neg_2av_1_22_port, neg_2a(21) => 
                           neg_2av_1_21_port, neg_2a(20) => neg_2av_1_20_port, 
                           neg_2a(19) => neg_2av_1_19_port, neg_2a(18) => 
                           neg_2av_1_18_port, neg_2a(17) => neg_2av_1_17_port, 
                           neg_2a(16) => neg_2av_1_16_port, neg_2a(15) => 
                           neg_2av_1_15_port, neg_2a(14) => neg_2av_1_14_port, 
                           neg_2a(13) => neg_2av_1_13_port, neg_2a(12) => 
                           neg_2av_1_12_port, neg_2a(11) => neg_2av_1_11_port, 
                           neg_2a(10) => neg_2av_1_10_port, neg_2a(9) => 
                           neg_2av_1_9_port, neg_2a(8) => neg_2av_1_8_port, 
                           neg_2a(7) => neg_2av_1_7_port, neg_2a(6) => 
                           neg_2av_1_6_port, neg_2a(5) => neg_2av_1_5_port, 
                           neg_2a(4) => neg_2av_1_4_port, neg_2a(3) => 
                           neg_2av_1_3_port, neg_2a(2) => neg_2av_1_2_port, 
                           neg_2a(1) => neg_2av_1_1_port, neg_2a(0) => 
                           neg_2av_1_0_port, sel(2) => b(3), sel(1) => b(2), 
                           sel(0) => b(1), s_out(31) => sum_vector_1_31_port, 
                           s_out(30) => sum_vector_1_30_port, s_out(29) => 
                           sum_vector_1_29_port, s_out(28) => 
                           sum_vector_1_28_port, s_out(27) => 
                           sum_vector_1_27_port, s_out(26) => 
                           sum_vector_1_26_port, s_out(25) => 
                           sum_vector_1_25_port, s_out(24) => 
                           sum_vector_1_24_port, s_out(23) => 
                           sum_vector_1_23_port, s_out(22) => 
                           sum_vector_1_22_port, s_out(21) => 
                           sum_vector_1_21_port, s_out(20) => 
                           sum_vector_1_20_port, s_out(19) => 
                           sum_vector_1_19_port, s_out(18) => 
                           sum_vector_1_18_port, s_out(17) => 
                           sum_vector_1_17_port, s_out(16) => 
                           sum_vector_1_16_port, s_out(15) => 
                           sum_vector_1_15_port, s_out(14) => 
                           sum_vector_1_14_port, s_out(13) => 
                           sum_vector_1_13_port, s_out(12) => 
                           sum_vector_1_12_port, s_out(11) => 
                           sum_vector_1_11_port, s_out(10) => 
                           sum_vector_1_10_port, s_out(9) => 
                           sum_vector_1_9_port, s_out(8) => sum_vector_1_8_port
                           , s_out(7) => sum_vector_1_7_port, s_out(6) => 
                           sum_vector_1_6_port, s_out(5) => sum_vector_1_5_port
                           , s_out(4) => sum_vector_1_4_port, s_out(3) => 
                           sum_vector_1_3_port, s_out(2) => sum_vector_1_2_port
                           , s_out(1) => sum_vector_1_1_port, s_out(0) => 
                           sum_vector_1_0_port);
   sum0_1 : rca_signed_NBIT32_0 port map( a(31) => sum_vector_0_31_port, a(30) 
                           => sum_vector_0_30_port, a(29) => 
                           sum_vector_0_29_port, a(28) => sum_vector_0_28_port,
                           a(27) => sum_vector_0_27_port, a(26) => 
                           sum_vector_0_26_port, a(25) => sum_vector_0_25_port,
                           a(24) => sum_vector_0_24_port, a(23) => 
                           sum_vector_0_23_port, a(22) => sum_vector_0_22_port,
                           a(21) => sum_vector_0_21_port, a(20) => 
                           sum_vector_0_20_port, a(19) => sum_vector_0_19_port,
                           a(18) => sum_vector_0_18_port, a(17) => 
                           sum_vector_0_17_port, a(16) => sum_vector_0_16_port,
                           a(15) => sum_vector_0_15_port, a(14) => 
                           sum_vector_0_14_port, a(13) => sum_vector_0_13_port,
                           a(12) => sum_vector_0_12_port, a(11) => 
                           sum_vector_0_11_port, a(10) => sum_vector_0_10_port,
                           a(9) => sum_vector_0_9_port, a(8) => 
                           sum_vector_0_8_port, a(7) => sum_vector_0_7_port, 
                           a(6) => sum_vector_0_6_port, a(5) => 
                           sum_vector_0_5_port, a(4) => sum_vector_0_4_port, 
                           a(3) => sum_vector_0_3_port, a(2) => 
                           sum_vector_0_2_port, a(1) => sum_vector_0_1_port, 
                           a(0) => sum_vector_0_0_port, b(31) => 
                           sum_vector_1_31_port, b(30) => sum_vector_1_30_port,
                           b(29) => sum_vector_1_29_port, b(28) => 
                           sum_vector_1_28_port, b(27) => sum_vector_1_27_port,
                           b(26) => sum_vector_1_26_port, b(25) => 
                           sum_vector_1_25_port, b(24) => sum_vector_1_24_port,
                           b(23) => sum_vector_1_23_port, b(22) => 
                           sum_vector_1_22_port, b(21) => sum_vector_1_21_port,
                           b(20) => sum_vector_1_20_port, b(19) => 
                           sum_vector_1_19_port, b(18) => sum_vector_1_18_port,
                           b(17) => sum_vector_1_17_port, b(16) => 
                           sum_vector_1_16_port, b(15) => sum_vector_1_15_port,
                           b(14) => sum_vector_1_14_port, b(13) => 
                           sum_vector_1_13_port, b(12) => sum_vector_1_12_port,
                           b(11) => sum_vector_1_11_port, b(10) => 
                           sum_vector_1_10_port, b(9) => sum_vector_1_9_port, 
                           b(8) => sum_vector_1_8_port, b(7) => 
                           sum_vector_1_7_port, b(6) => sum_vector_1_6_port, 
                           b(5) => sum_vector_1_5_port, b(4) => 
                           sum_vector_1_4_port, b(3) => sum_vector_1_3_port, 
                           b(2) => sum_vector_1_2_port, b(1) => 
                           sum_vector_1_1_port, b(0) => sum_vector_1_0_port, c 
                           => n_1176, s(31) => sum_vector_2_31_port, s(30) => 
                           sum_vector_2_30_port, s(29) => sum_vector_2_29_port,
                           s(28) => sum_vector_2_28_port, s(27) => 
                           sum_vector_2_27_port, s(26) => sum_vector_2_26_port,
                           s(25) => sum_vector_2_25_port, s(24) => 
                           sum_vector_2_24_port, s(23) => sum_vector_2_23_port,
                           s(22) => sum_vector_2_22_port, s(21) => 
                           sum_vector_2_21_port, s(20) => sum_vector_2_20_port,
                           s(19) => sum_vector_2_19_port, s(18) => 
                           sum_vector_2_18_port, s(17) => sum_vector_2_17_port,
                           s(16) => sum_vector_2_16_port, s(15) => 
                           sum_vector_2_15_port, s(14) => sum_vector_2_14_port,
                           s(13) => sum_vector_2_13_port, s(12) => 
                           sum_vector_2_12_port, s(11) => sum_vector_2_11_port,
                           s(10) => sum_vector_2_10_port, s(9) => 
                           sum_vector_2_9_port, s(8) => sum_vector_2_8_port, 
                           s(7) => sum_vector_2_7_port, s(6) => 
                           sum_vector_2_6_port, s(5) => sum_vector_2_5_port, 
                           s(4) => sum_vector_2_4_port, s(3) => 
                           sum_vector_2_3_port, s(2) => sum_vector_2_2_port, 
                           s(1) => sum_vector_2_1_port, s(0) => 
                           sum_vector_2_0_port);
   shn_2 : shift_NBIT32_SHIFT2 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_2_31_port, pos_a(30) => 
                           pos_av_2_30_port, pos_a(29) => pos_av_2_29_port, 
                           pos_a(28) => pos_av_2_28_port, pos_a(27) => 
                           pos_av_2_27_port, pos_a(26) => pos_av_2_26_port, 
                           pos_a(25) => pos_av_2_25_port, pos_a(24) => 
                           pos_av_2_24_port, pos_a(23) => pos_av_2_23_port, 
                           pos_a(22) => pos_av_2_22_port, pos_a(21) => 
                           pos_av_2_21_port, pos_a(20) => pos_av_2_20_port, 
                           pos_a(19) => pos_av_2_19_port, pos_a(18) => 
                           pos_av_2_18_port, pos_a(17) => pos_av_2_17_port, 
                           pos_a(16) => pos_av_2_16_port, pos_a(15) => 
                           pos_av_2_15_port, pos_a(14) => pos_av_2_14_port, 
                           pos_a(13) => pos_av_2_13_port, pos_a(12) => 
                           pos_av_2_12_port, pos_a(11) => pos_av_2_11_port, 
                           pos_a(10) => pos_av_2_10_port, pos_a(9) => 
                           pos_av_2_9_port, pos_a(8) => pos_av_2_8_port, 
                           pos_a(7) => pos_av_2_7_port, pos_a(6) => 
                           pos_av_2_6_port, pos_a(5) => pos_av_2_5_port, 
                           pos_a(4) => pos_av_2_4_port, pos_a(3) => n_1177, 
                           pos_a(2) => n_1178, pos_a(1) => n_1179, pos_a(0) => 
                           n_1180, neg_a(31) => neg_av_2_31_port, neg_a(30) => 
                           neg_av_2_30_port, neg_a(29) => neg_av_2_29_port, 
                           neg_a(28) => neg_av_2_28_port, neg_a(27) => 
                           neg_av_2_27_port, neg_a(26) => neg_av_2_26_port, 
                           neg_a(25) => neg_av_2_25_port, neg_a(24) => 
                           neg_av_2_24_port, neg_a(23) => neg_av_2_23_port, 
                           neg_a(22) => neg_av_2_22_port, neg_a(21) => 
                           neg_av_2_21_port, neg_a(20) => neg_av_2_20_port, 
                           neg_a(19) => neg_av_2_19_port, neg_a(18) => 
                           neg_av_2_18_port, neg_a(17) => neg_av_2_17_port, 
                           neg_a(16) => neg_av_2_16_port, neg_a(15) => 
                           neg_av_2_15_port, neg_a(14) => neg_av_2_14_port, 
                           neg_a(13) => neg_av_2_13_port, neg_a(12) => 
                           neg_av_2_12_port, neg_a(11) => neg_av_2_11_port, 
                           neg_a(10) => neg_av_2_10_port, neg_a(9) => 
                           neg_av_2_9_port, neg_a(8) => neg_av_2_8_port, 
                           neg_a(7) => neg_av_2_7_port, neg_a(6) => 
                           neg_av_2_6_port, neg_a(5) => neg_av_2_5_port, 
                           neg_a(4) => neg_av_2_4_port, neg_a(3) => n_1181, 
                           neg_a(2) => n_1182, neg_a(1) => n_1183, neg_a(0) => 
                           n_1184, pos_2a(31) => pos_2av_2_31_port, pos_2a(30) 
                           => pos_2av_2_30_port, pos_2a(29) => 
                           pos_2av_2_29_port, pos_2a(28) => pos_2av_2_28_port, 
                           pos_2a(27) => pos_2av_2_27_port, pos_2a(26) => 
                           pos_2av_2_26_port, pos_2a(25) => pos_2av_2_25_port, 
                           pos_2a(24) => pos_2av_2_24_port, pos_2a(23) => 
                           pos_2av_2_23_port, pos_2a(22) => pos_2av_2_22_port, 
                           pos_2a(21) => pos_2av_2_21_port, pos_2a(20) => 
                           pos_2av_2_20_port, pos_2a(19) => pos_2av_2_19_port, 
                           pos_2a(18) => pos_2av_2_18_port, pos_2a(17) => 
                           pos_2av_2_17_port, pos_2a(16) => pos_2av_2_16_port, 
                           pos_2a(15) => pos_2av_2_15_port, pos_2a(14) => 
                           pos_2av_2_14_port, pos_2a(13) => pos_2av_2_13_port, 
                           pos_2a(12) => pos_2av_2_12_port, pos_2a(11) => 
                           pos_2av_2_11_port, pos_2a(10) => pos_2av_2_10_port, 
                           pos_2a(9) => pos_2av_2_9_port, pos_2a(8) => 
                           pos_2av_2_8_port, pos_2a(7) => pos_2av_2_7_port, 
                           pos_2a(6) => pos_2av_2_6_port, pos_2a(5) => 
                           pos_2av_2_5_port, pos_2a(4) => n_1185, pos_2a(3) => 
                           n_1186, pos_2a(2) => n_1187, pos_2a(1) => n_1188, 
                           pos_2a(0) => n_1189, neg_2a(31) => neg_2av_2_31_port
                           , neg_2a(30) => neg_2av_2_30_port, neg_2a(29) => 
                           neg_2av_2_29_port, neg_2a(28) => neg_2av_2_28_port, 
                           neg_2a(27) => neg_2av_2_27_port, neg_2a(26) => 
                           neg_2av_2_26_port, neg_2a(25) => neg_2av_2_25_port, 
                           neg_2a(24) => neg_2av_2_24_port, neg_2a(23) => 
                           neg_2av_2_23_port, neg_2a(22) => neg_2av_2_22_port, 
                           neg_2a(21) => neg_2av_2_21_port, neg_2a(20) => 
                           neg_2av_2_20_port, neg_2a(19) => neg_2av_2_19_port, 
                           neg_2a(18) => neg_2av_2_18_port, neg_2a(17) => 
                           neg_2av_2_17_port, neg_2a(16) => neg_2av_2_16_port, 
                           neg_2a(15) => neg_2av_2_15_port, neg_2a(14) => 
                           neg_2av_2_14_port, neg_2a(13) => neg_2av_2_13_port, 
                           neg_2a(12) => neg_2av_2_12_port, neg_2a(11) => 
                           neg_2av_2_11_port, neg_2a(10) => neg_2av_2_10_port, 
                           neg_2a(9) => neg_2av_2_9_port, neg_2a(8) => 
                           neg_2av_2_8_port, neg_2a(7) => neg_2av_2_7_port, 
                           neg_2a(6) => neg_2av_2_6_port, neg_2a(5) => 
                           neg_2av_2_5_port, neg_2a(4) => n_1190, neg_2a(3) => 
                           n_1191, neg_2a(2) => n_1192, neg_2a(1) => n_1193, 
                           neg_2a(0) => n_1194);
   vpn_2 : vp_NBIT32_6 port map( pos_a(31) => pos_av_2_31_port, pos_a(30) => 
                           pos_av_2_30_port, pos_a(29) => pos_av_2_29_port, 
                           pos_a(28) => pos_av_2_28_port, pos_a(27) => 
                           pos_av_2_27_port, pos_a(26) => pos_av_2_26_port, 
                           pos_a(25) => pos_av_2_25_port, pos_a(24) => 
                           pos_av_2_24_port, pos_a(23) => pos_av_2_23_port, 
                           pos_a(22) => pos_av_2_22_port, pos_a(21) => 
                           pos_av_2_21_port, pos_a(20) => pos_av_2_20_port, 
                           pos_a(19) => pos_av_2_19_port, pos_a(18) => 
                           pos_av_2_18_port, pos_a(17) => pos_av_2_17_port, 
                           pos_a(16) => pos_av_2_16_port, pos_a(15) => 
                           pos_av_2_15_port, pos_a(14) => pos_av_2_14_port, 
                           pos_a(13) => pos_av_2_13_port, pos_a(12) => 
                           pos_av_2_12_port, pos_a(11) => pos_av_2_11_port, 
                           pos_a(10) => pos_av_2_10_port, pos_a(9) => 
                           pos_av_2_9_port, pos_a(8) => pos_av_2_8_port, 
                           pos_a(7) => pos_av_2_7_port, pos_a(6) => 
                           pos_av_2_6_port, pos_a(5) => pos_av_2_5_port, 
                           pos_a(4) => pos_av_2_4_port, pos_a(3) => 
                           pos_av_2_3_port, pos_a(2) => pos_av_2_2_port, 
                           pos_a(1) => pos_av_2_1_port, pos_a(0) => 
                           pos_av_2_0_port, neg_a(31) => neg_av_2_31_port, 
                           neg_a(30) => neg_av_2_30_port, neg_a(29) => 
                           neg_av_2_29_port, neg_a(28) => neg_av_2_28_port, 
                           neg_a(27) => neg_av_2_27_port, neg_a(26) => 
                           neg_av_2_26_port, neg_a(25) => neg_av_2_25_port, 
                           neg_a(24) => neg_av_2_24_port, neg_a(23) => 
                           neg_av_2_23_port, neg_a(22) => neg_av_2_22_port, 
                           neg_a(21) => neg_av_2_21_port, neg_a(20) => 
                           neg_av_2_20_port, neg_a(19) => neg_av_2_19_port, 
                           neg_a(18) => neg_av_2_18_port, neg_a(17) => 
                           neg_av_2_17_port, neg_a(16) => neg_av_2_16_port, 
                           neg_a(15) => neg_av_2_15_port, neg_a(14) => 
                           neg_av_2_14_port, neg_a(13) => neg_av_2_13_port, 
                           neg_a(12) => neg_av_2_12_port, neg_a(11) => 
                           neg_av_2_11_port, neg_a(10) => neg_av_2_10_port, 
                           neg_a(9) => neg_av_2_9_port, neg_a(8) => 
                           neg_av_2_8_port, neg_a(7) => neg_av_2_7_port, 
                           neg_a(6) => neg_av_2_6_port, neg_a(5) => 
                           neg_av_2_5_port, neg_a(4) => neg_av_2_4_port, 
                           neg_a(3) => neg_av_2_3_port, neg_a(2) => 
                           neg_av_2_2_port, neg_a(1) => neg_av_2_1_port, 
                           neg_a(0) => neg_av_2_0_port, pos_2a(31) => 
                           pos_2av_2_31_port, pos_2a(30) => pos_2av_2_30_port, 
                           pos_2a(29) => pos_2av_2_29_port, pos_2a(28) => 
                           pos_2av_2_28_port, pos_2a(27) => pos_2av_2_27_port, 
                           pos_2a(26) => pos_2av_2_26_port, pos_2a(25) => 
                           pos_2av_2_25_port, pos_2a(24) => pos_2av_2_24_port, 
                           pos_2a(23) => pos_2av_2_23_port, pos_2a(22) => 
                           pos_2av_2_22_port, pos_2a(21) => pos_2av_2_21_port, 
                           pos_2a(20) => pos_2av_2_20_port, pos_2a(19) => 
                           pos_2av_2_19_port, pos_2a(18) => pos_2av_2_18_port, 
                           pos_2a(17) => pos_2av_2_17_port, pos_2a(16) => 
                           pos_2av_2_16_port, pos_2a(15) => pos_2av_2_15_port, 
                           pos_2a(14) => pos_2av_2_14_port, pos_2a(13) => 
                           pos_2av_2_13_port, pos_2a(12) => pos_2av_2_12_port, 
                           pos_2a(11) => pos_2av_2_11_port, pos_2a(10) => 
                           pos_2av_2_10_port, pos_2a(9) => pos_2av_2_9_port, 
                           pos_2a(8) => pos_2av_2_8_port, pos_2a(7) => 
                           pos_2av_2_7_port, pos_2a(6) => pos_2av_2_6_port, 
                           pos_2a(5) => pos_2av_2_5_port, pos_2a(4) => 
                           pos_2av_2_4_port, pos_2a(3) => pos_2av_2_3_port, 
                           pos_2a(2) => pos_2av_2_2_port, pos_2a(1) => 
                           pos_2av_2_1_port, pos_2a(0) => pos_2av_2_0_port, 
                           neg_2a(31) => neg_2av_2_31_port, neg_2a(30) => 
                           neg_2av_2_30_port, neg_2a(29) => neg_2av_2_29_port, 
                           neg_2a(28) => neg_2av_2_28_port, neg_2a(27) => 
                           neg_2av_2_27_port, neg_2a(26) => neg_2av_2_26_port, 
                           neg_2a(25) => neg_2av_2_25_port, neg_2a(24) => 
                           neg_2av_2_24_port, neg_2a(23) => neg_2av_2_23_port, 
                           neg_2a(22) => neg_2av_2_22_port, neg_2a(21) => 
                           neg_2av_2_21_port, neg_2a(20) => neg_2av_2_20_port, 
                           neg_2a(19) => neg_2av_2_19_port, neg_2a(18) => 
                           neg_2av_2_18_port, neg_2a(17) => neg_2av_2_17_port, 
                           neg_2a(16) => neg_2av_2_16_port, neg_2a(15) => 
                           neg_2av_2_15_port, neg_2a(14) => neg_2av_2_14_port, 
                           neg_2a(13) => neg_2av_2_13_port, neg_2a(12) => 
                           neg_2av_2_12_port, neg_2a(11) => neg_2av_2_11_port, 
                           neg_2a(10) => neg_2av_2_10_port, neg_2a(9) => 
                           neg_2av_2_9_port, neg_2a(8) => neg_2av_2_8_port, 
                           neg_2a(7) => neg_2av_2_7_port, neg_2a(6) => 
                           neg_2av_2_6_port, neg_2a(5) => neg_2av_2_5_port, 
                           neg_2a(4) => neg_2av_2_4_port, neg_2a(3) => 
                           neg_2av_2_3_port, neg_2a(2) => neg_2av_2_2_port, 
                           neg_2a(1) => neg_2av_2_1_port, neg_2a(0) => 
                           neg_2av_2_0_port, sel(2) => b(5), sel(1) => b(4), 
                           sel(0) => b(3), s_out(31) => sum_vector_3_31_port, 
                           s_out(30) => sum_vector_3_30_port, s_out(29) => 
                           sum_vector_3_29_port, s_out(28) => 
                           sum_vector_3_28_port, s_out(27) => 
                           sum_vector_3_27_port, s_out(26) => 
                           sum_vector_3_26_port, s_out(25) => 
                           sum_vector_3_25_port, s_out(24) => 
                           sum_vector_3_24_port, s_out(23) => 
                           sum_vector_3_23_port, s_out(22) => 
                           sum_vector_3_22_port, s_out(21) => 
                           sum_vector_3_21_port, s_out(20) => 
                           sum_vector_3_20_port, s_out(19) => 
                           sum_vector_3_19_port, s_out(18) => 
                           sum_vector_3_18_port, s_out(17) => 
                           sum_vector_3_17_port, s_out(16) => 
                           sum_vector_3_16_port, s_out(15) => 
                           sum_vector_3_15_port, s_out(14) => 
                           sum_vector_3_14_port, s_out(13) => 
                           sum_vector_3_13_port, s_out(12) => 
                           sum_vector_3_12_port, s_out(11) => 
                           sum_vector_3_11_port, s_out(10) => 
                           sum_vector_3_10_port, s_out(9) => 
                           sum_vector_3_9_port, s_out(8) => sum_vector_3_8_port
                           , s_out(7) => sum_vector_3_7_port, s_out(6) => 
                           sum_vector_3_6_port, s_out(5) => sum_vector_3_5_port
                           , s_out(4) => sum_vector_3_4_port, s_out(3) => 
                           sum_vector_3_3_port, s_out(2) => sum_vector_3_2_port
                           , s_out(1) => sum_vector_3_1_port, s_out(0) => 
                           sum_vector_3_0_port);
   sumn_2 : rca_signed_NBIT32_6 port map( a(31) => sum_vector_2_31_port, a(30) 
                           => sum_vector_2_30_port, a(29) => 
                           sum_vector_2_29_port, a(28) => sum_vector_2_28_port,
                           a(27) => sum_vector_2_27_port, a(26) => 
                           sum_vector_2_26_port, a(25) => sum_vector_2_25_port,
                           a(24) => sum_vector_2_24_port, a(23) => 
                           sum_vector_2_23_port, a(22) => sum_vector_2_22_port,
                           a(21) => sum_vector_2_21_port, a(20) => 
                           sum_vector_2_20_port, a(19) => sum_vector_2_19_port,
                           a(18) => sum_vector_2_18_port, a(17) => 
                           sum_vector_2_17_port, a(16) => sum_vector_2_16_port,
                           a(15) => sum_vector_2_15_port, a(14) => 
                           sum_vector_2_14_port, a(13) => sum_vector_2_13_port,
                           a(12) => sum_vector_2_12_port, a(11) => 
                           sum_vector_2_11_port, a(10) => sum_vector_2_10_port,
                           a(9) => sum_vector_2_9_port, a(8) => 
                           sum_vector_2_8_port, a(7) => sum_vector_2_7_port, 
                           a(6) => sum_vector_2_6_port, a(5) => 
                           sum_vector_2_5_port, a(4) => sum_vector_2_4_port, 
                           a(3) => sum_vector_2_3_port, a(2) => 
                           sum_vector_2_2_port, a(1) => sum_vector_2_1_port, 
                           a(0) => sum_vector_2_0_port, b(31) => 
                           sum_vector_3_31_port, b(30) => sum_vector_3_30_port,
                           b(29) => sum_vector_3_29_port, b(28) => 
                           sum_vector_3_28_port, b(27) => sum_vector_3_27_port,
                           b(26) => sum_vector_3_26_port, b(25) => 
                           sum_vector_3_25_port, b(24) => sum_vector_3_24_port,
                           b(23) => sum_vector_3_23_port, b(22) => 
                           sum_vector_3_22_port, b(21) => sum_vector_3_21_port,
                           b(20) => sum_vector_3_20_port, b(19) => 
                           sum_vector_3_19_port, b(18) => sum_vector_3_18_port,
                           b(17) => sum_vector_3_17_port, b(16) => 
                           sum_vector_3_16_port, b(15) => sum_vector_3_15_port,
                           b(14) => sum_vector_3_14_port, b(13) => 
                           sum_vector_3_13_port, b(12) => sum_vector_3_12_port,
                           b(11) => sum_vector_3_11_port, b(10) => 
                           sum_vector_3_10_port, b(9) => sum_vector_3_9_port, 
                           b(8) => sum_vector_3_8_port, b(7) => 
                           sum_vector_3_7_port, b(6) => sum_vector_3_6_port, 
                           b(5) => sum_vector_3_5_port, b(4) => 
                           sum_vector_3_4_port, b(3) => sum_vector_3_3_port, 
                           b(2) => sum_vector_3_2_port, b(1) => 
                           sum_vector_3_1_port, b(0) => sum_vector_3_0_port, c 
                           => n_1195, s(31) => sum_vector_4_31_port, s(30) => 
                           sum_vector_4_30_port, s(29) => sum_vector_4_29_port,
                           s(28) => sum_vector_4_28_port, s(27) => 
                           sum_vector_4_27_port, s(26) => sum_vector_4_26_port,
                           s(25) => sum_vector_4_25_port, s(24) => 
                           sum_vector_4_24_port, s(23) => sum_vector_4_23_port,
                           s(22) => sum_vector_4_22_port, s(21) => 
                           sum_vector_4_21_port, s(20) => sum_vector_4_20_port,
                           s(19) => sum_vector_4_19_port, s(18) => 
                           sum_vector_4_18_port, s(17) => sum_vector_4_17_port,
                           s(16) => sum_vector_4_16_port, s(15) => 
                           sum_vector_4_15_port, s(14) => sum_vector_4_14_port,
                           s(13) => sum_vector_4_13_port, s(12) => 
                           sum_vector_4_12_port, s(11) => sum_vector_4_11_port,
                           s(10) => sum_vector_4_10_port, s(9) => 
                           sum_vector_4_9_port, s(8) => sum_vector_4_8_port, 
                           s(7) => sum_vector_4_7_port, s(6) => 
                           sum_vector_4_6_port, s(5) => sum_vector_4_5_port, 
                           s(4) => sum_vector_4_4_port, s(3) => 
                           sum_vector_4_3_port, s(2) => sum_vector_4_2_port, 
                           s(1) => sum_vector_4_1_port, s(0) => 
                           sum_vector_4_0_port);
   shn_3 : shift_NBIT32_SHIFT3 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_3_31_port, pos_a(30) => 
                           pos_av_3_30_port, pos_a(29) => pos_av_3_29_port, 
                           pos_a(28) => pos_av_3_28_port, pos_a(27) => 
                           pos_av_3_27_port, pos_a(26) => pos_av_3_26_port, 
                           pos_a(25) => pos_av_3_25_port, pos_a(24) => 
                           pos_av_3_24_port, pos_a(23) => pos_av_3_23_port, 
                           pos_a(22) => pos_av_3_22_port, pos_a(21) => 
                           pos_av_3_21_port, pos_a(20) => pos_av_3_20_port, 
                           pos_a(19) => pos_av_3_19_port, pos_a(18) => 
                           pos_av_3_18_port, pos_a(17) => pos_av_3_17_port, 
                           pos_a(16) => pos_av_3_16_port, pos_a(15) => 
                           pos_av_3_15_port, pos_a(14) => pos_av_3_14_port, 
                           pos_a(13) => pos_av_3_13_port, pos_a(12) => 
                           pos_av_3_12_port, pos_a(11) => pos_av_3_11_port, 
                           pos_a(10) => pos_av_3_10_port, pos_a(9) => 
                           pos_av_3_9_port, pos_a(8) => pos_av_3_8_port, 
                           pos_a(7) => pos_av_3_7_port, pos_a(6) => 
                           pos_av_3_6_port, pos_a(5) => n_1196, pos_a(4) => 
                           n_1197, pos_a(3) => n_1198, pos_a(2) => n_1199, 
                           pos_a(1) => n_1200, pos_a(0) => n_1201, neg_a(31) =>
                           neg_av_3_31_port, neg_a(30) => neg_av_3_30_port, 
                           neg_a(29) => neg_av_3_29_port, neg_a(28) => 
                           neg_av_3_28_port, neg_a(27) => neg_av_3_27_port, 
                           neg_a(26) => neg_av_3_26_port, neg_a(25) => 
                           neg_av_3_25_port, neg_a(24) => neg_av_3_24_port, 
                           neg_a(23) => neg_av_3_23_port, neg_a(22) => 
                           neg_av_3_22_port, neg_a(21) => neg_av_3_21_port, 
                           neg_a(20) => neg_av_3_20_port, neg_a(19) => 
                           neg_av_3_19_port, neg_a(18) => neg_av_3_18_port, 
                           neg_a(17) => neg_av_3_17_port, neg_a(16) => 
                           neg_av_3_16_port, neg_a(15) => neg_av_3_15_port, 
                           neg_a(14) => neg_av_3_14_port, neg_a(13) => 
                           neg_av_3_13_port, neg_a(12) => neg_av_3_12_port, 
                           neg_a(11) => neg_av_3_11_port, neg_a(10) => 
                           neg_av_3_10_port, neg_a(9) => neg_av_3_9_port, 
                           neg_a(8) => neg_av_3_8_port, neg_a(7) => 
                           neg_av_3_7_port, neg_a(6) => neg_av_3_6_port, 
                           neg_a(5) => n_1202, neg_a(4) => n_1203, neg_a(3) => 
                           n_1204, neg_a(2) => n_1205, neg_a(1) => n_1206, 
                           neg_a(0) => n_1207, pos_2a(31) => pos_2av_3_31_port,
                           pos_2a(30) => pos_2av_3_30_port, pos_2a(29) => 
                           pos_2av_3_29_port, pos_2a(28) => pos_2av_3_28_port, 
                           pos_2a(27) => pos_2av_3_27_port, pos_2a(26) => 
                           pos_2av_3_26_port, pos_2a(25) => pos_2av_3_25_port, 
                           pos_2a(24) => pos_2av_3_24_port, pos_2a(23) => 
                           pos_2av_3_23_port, pos_2a(22) => pos_2av_3_22_port, 
                           pos_2a(21) => pos_2av_3_21_port, pos_2a(20) => 
                           pos_2av_3_20_port, pos_2a(19) => pos_2av_3_19_port, 
                           pos_2a(18) => pos_2av_3_18_port, pos_2a(17) => 
                           pos_2av_3_17_port, pos_2a(16) => pos_2av_3_16_port, 
                           pos_2a(15) => pos_2av_3_15_port, pos_2a(14) => 
                           pos_2av_3_14_port, pos_2a(13) => pos_2av_3_13_port, 
                           pos_2a(12) => pos_2av_3_12_port, pos_2a(11) => 
                           pos_2av_3_11_port, pos_2a(10) => pos_2av_3_10_port, 
                           pos_2a(9) => pos_2av_3_9_port, pos_2a(8) => 
                           pos_2av_3_8_port, pos_2a(7) => pos_2av_3_7_port, 
                           pos_2a(6) => n_1208, pos_2a(5) => n_1209, pos_2a(4) 
                           => n_1210, pos_2a(3) => n_1211, pos_2a(2) => n_1212,
                           pos_2a(1) => n_1213, pos_2a(0) => n_1214, neg_2a(31)
                           => neg_2av_3_31_port, neg_2a(30) => 
                           neg_2av_3_30_port, neg_2a(29) => neg_2av_3_29_port, 
                           neg_2a(28) => neg_2av_3_28_port, neg_2a(27) => 
                           neg_2av_3_27_port, neg_2a(26) => neg_2av_3_26_port, 
                           neg_2a(25) => neg_2av_3_25_port, neg_2a(24) => 
                           neg_2av_3_24_port, neg_2a(23) => neg_2av_3_23_port, 
                           neg_2a(22) => neg_2av_3_22_port, neg_2a(21) => 
                           neg_2av_3_21_port, neg_2a(20) => neg_2av_3_20_port, 
                           neg_2a(19) => neg_2av_3_19_port, neg_2a(18) => 
                           neg_2av_3_18_port, neg_2a(17) => neg_2av_3_17_port, 
                           neg_2a(16) => neg_2av_3_16_port, neg_2a(15) => 
                           neg_2av_3_15_port, neg_2a(14) => neg_2av_3_14_port, 
                           neg_2a(13) => neg_2av_3_13_port, neg_2a(12) => 
                           neg_2av_3_12_port, neg_2a(11) => neg_2av_3_11_port, 
                           neg_2a(10) => neg_2av_3_10_port, neg_2a(9) => 
                           neg_2av_3_9_port, neg_2a(8) => neg_2av_3_8_port, 
                           neg_2a(7) => neg_2av_3_7_port, neg_2a(6) => n_1215, 
                           neg_2a(5) => n_1216, neg_2a(4) => n_1217, neg_2a(3) 
                           => n_1218, neg_2a(2) => n_1219, neg_2a(1) => n_1220,
                           neg_2a(0) => n_1221);
   vpn_3 : vp_NBIT32_5 port map( pos_a(31) => pos_av_3_31_port, pos_a(30) => 
                           pos_av_3_30_port, pos_a(29) => pos_av_3_29_port, 
                           pos_a(28) => pos_av_3_28_port, pos_a(27) => 
                           pos_av_3_27_port, pos_a(26) => pos_av_3_26_port, 
                           pos_a(25) => pos_av_3_25_port, pos_a(24) => 
                           pos_av_3_24_port, pos_a(23) => pos_av_3_23_port, 
                           pos_a(22) => pos_av_3_22_port, pos_a(21) => 
                           pos_av_3_21_port, pos_a(20) => pos_av_3_20_port, 
                           pos_a(19) => pos_av_3_19_port, pos_a(18) => 
                           pos_av_3_18_port, pos_a(17) => pos_av_3_17_port, 
                           pos_a(16) => pos_av_3_16_port, pos_a(15) => 
                           pos_av_3_15_port, pos_a(14) => pos_av_3_14_port, 
                           pos_a(13) => pos_av_3_13_port, pos_a(12) => 
                           pos_av_3_12_port, pos_a(11) => pos_av_3_11_port, 
                           pos_a(10) => pos_av_3_10_port, pos_a(9) => 
                           pos_av_3_9_port, pos_a(8) => pos_av_3_8_port, 
                           pos_a(7) => pos_av_3_7_port, pos_a(6) => 
                           pos_av_3_6_port, pos_a(5) => pos_av_3_5_port, 
                           pos_a(4) => pos_av_3_4_port, pos_a(3) => 
                           pos_av_3_3_port, pos_a(2) => pos_av_3_2_port, 
                           pos_a(1) => pos_av_3_1_port, pos_a(0) => 
                           pos_av_3_0_port, neg_a(31) => neg_av_3_31_port, 
                           neg_a(30) => neg_av_3_30_port, neg_a(29) => 
                           neg_av_3_29_port, neg_a(28) => neg_av_3_28_port, 
                           neg_a(27) => neg_av_3_27_port, neg_a(26) => 
                           neg_av_3_26_port, neg_a(25) => neg_av_3_25_port, 
                           neg_a(24) => neg_av_3_24_port, neg_a(23) => 
                           neg_av_3_23_port, neg_a(22) => neg_av_3_22_port, 
                           neg_a(21) => neg_av_3_21_port, neg_a(20) => 
                           neg_av_3_20_port, neg_a(19) => neg_av_3_19_port, 
                           neg_a(18) => neg_av_3_18_port, neg_a(17) => 
                           neg_av_3_17_port, neg_a(16) => neg_av_3_16_port, 
                           neg_a(15) => neg_av_3_15_port, neg_a(14) => 
                           neg_av_3_14_port, neg_a(13) => neg_av_3_13_port, 
                           neg_a(12) => neg_av_3_12_port, neg_a(11) => 
                           neg_av_3_11_port, neg_a(10) => neg_av_3_10_port, 
                           neg_a(9) => neg_av_3_9_port, neg_a(8) => 
                           neg_av_3_8_port, neg_a(7) => neg_av_3_7_port, 
                           neg_a(6) => neg_av_3_6_port, neg_a(5) => 
                           neg_av_3_5_port, neg_a(4) => neg_av_3_4_port, 
                           neg_a(3) => neg_av_3_3_port, neg_a(2) => 
                           neg_av_3_2_port, neg_a(1) => neg_av_3_1_port, 
                           neg_a(0) => neg_av_3_0_port, pos_2a(31) => 
                           pos_2av_3_31_port, pos_2a(30) => pos_2av_3_30_port, 
                           pos_2a(29) => pos_2av_3_29_port, pos_2a(28) => 
                           pos_2av_3_28_port, pos_2a(27) => pos_2av_3_27_port, 
                           pos_2a(26) => pos_2av_3_26_port, pos_2a(25) => 
                           pos_2av_3_25_port, pos_2a(24) => pos_2av_3_24_port, 
                           pos_2a(23) => pos_2av_3_23_port, pos_2a(22) => 
                           pos_2av_3_22_port, pos_2a(21) => pos_2av_3_21_port, 
                           pos_2a(20) => pos_2av_3_20_port, pos_2a(19) => 
                           pos_2av_3_19_port, pos_2a(18) => pos_2av_3_18_port, 
                           pos_2a(17) => pos_2av_3_17_port, pos_2a(16) => 
                           pos_2av_3_16_port, pos_2a(15) => pos_2av_3_15_port, 
                           pos_2a(14) => pos_2av_3_14_port, pos_2a(13) => 
                           pos_2av_3_13_port, pos_2a(12) => pos_2av_3_12_port, 
                           pos_2a(11) => pos_2av_3_11_port, pos_2a(10) => 
                           pos_2av_3_10_port, pos_2a(9) => pos_2av_3_9_port, 
                           pos_2a(8) => pos_2av_3_8_port, pos_2a(7) => 
                           pos_2av_3_7_port, pos_2a(6) => pos_2av_3_6_port, 
                           pos_2a(5) => pos_2av_3_5_port, pos_2a(4) => 
                           pos_2av_3_4_port, pos_2a(3) => pos_2av_3_3_port, 
                           pos_2a(2) => pos_2av_3_2_port, pos_2a(1) => 
                           pos_2av_3_1_port, pos_2a(0) => pos_2av_3_0_port, 
                           neg_2a(31) => neg_2av_3_31_port, neg_2a(30) => 
                           neg_2av_3_30_port, neg_2a(29) => neg_2av_3_29_port, 
                           neg_2a(28) => neg_2av_3_28_port, neg_2a(27) => 
                           neg_2av_3_27_port, neg_2a(26) => neg_2av_3_26_port, 
                           neg_2a(25) => neg_2av_3_25_port, neg_2a(24) => 
                           neg_2av_3_24_port, neg_2a(23) => neg_2av_3_23_port, 
                           neg_2a(22) => neg_2av_3_22_port, neg_2a(21) => 
                           neg_2av_3_21_port, neg_2a(20) => neg_2av_3_20_port, 
                           neg_2a(19) => neg_2av_3_19_port, neg_2a(18) => 
                           neg_2av_3_18_port, neg_2a(17) => neg_2av_3_17_port, 
                           neg_2a(16) => neg_2av_3_16_port, neg_2a(15) => 
                           neg_2av_3_15_port, neg_2a(14) => neg_2av_3_14_port, 
                           neg_2a(13) => neg_2av_3_13_port, neg_2a(12) => 
                           neg_2av_3_12_port, neg_2a(11) => neg_2av_3_11_port, 
                           neg_2a(10) => neg_2av_3_10_port, neg_2a(9) => 
                           neg_2av_3_9_port, neg_2a(8) => neg_2av_3_8_port, 
                           neg_2a(7) => neg_2av_3_7_port, neg_2a(6) => 
                           neg_2av_3_6_port, neg_2a(5) => neg_2av_3_5_port, 
                           neg_2a(4) => neg_2av_3_4_port, neg_2a(3) => 
                           neg_2av_3_3_port, neg_2a(2) => neg_2av_3_2_port, 
                           neg_2a(1) => neg_2av_3_1_port, neg_2a(0) => 
                           neg_2av_3_0_port, sel(2) => b(7), sel(1) => b(6), 
                           sel(0) => b(5), s_out(31) => sum_vector_5_31_port, 
                           s_out(30) => sum_vector_5_30_port, s_out(29) => 
                           sum_vector_5_29_port, s_out(28) => 
                           sum_vector_5_28_port, s_out(27) => 
                           sum_vector_5_27_port, s_out(26) => 
                           sum_vector_5_26_port, s_out(25) => 
                           sum_vector_5_25_port, s_out(24) => 
                           sum_vector_5_24_port, s_out(23) => 
                           sum_vector_5_23_port, s_out(22) => 
                           sum_vector_5_22_port, s_out(21) => 
                           sum_vector_5_21_port, s_out(20) => 
                           sum_vector_5_20_port, s_out(19) => 
                           sum_vector_5_19_port, s_out(18) => 
                           sum_vector_5_18_port, s_out(17) => 
                           sum_vector_5_17_port, s_out(16) => 
                           sum_vector_5_16_port, s_out(15) => 
                           sum_vector_5_15_port, s_out(14) => 
                           sum_vector_5_14_port, s_out(13) => 
                           sum_vector_5_13_port, s_out(12) => 
                           sum_vector_5_12_port, s_out(11) => 
                           sum_vector_5_11_port, s_out(10) => 
                           sum_vector_5_10_port, s_out(9) => 
                           sum_vector_5_9_port, s_out(8) => sum_vector_5_8_port
                           , s_out(7) => sum_vector_5_7_port, s_out(6) => 
                           sum_vector_5_6_port, s_out(5) => sum_vector_5_5_port
                           , s_out(4) => sum_vector_5_4_port, s_out(3) => 
                           sum_vector_5_3_port, s_out(2) => sum_vector_5_2_port
                           , s_out(1) => sum_vector_5_1_port, s_out(0) => 
                           sum_vector_5_0_port);
   sumn_3 : rca_signed_NBIT32_5 port map( a(31) => sum_vector_4_31_port, a(30) 
                           => sum_vector_4_30_port, a(29) => 
                           sum_vector_4_29_port, a(28) => sum_vector_4_28_port,
                           a(27) => sum_vector_4_27_port, a(26) => 
                           sum_vector_4_26_port, a(25) => sum_vector_4_25_port,
                           a(24) => sum_vector_4_24_port, a(23) => 
                           sum_vector_4_23_port, a(22) => sum_vector_4_22_port,
                           a(21) => sum_vector_4_21_port, a(20) => 
                           sum_vector_4_20_port, a(19) => sum_vector_4_19_port,
                           a(18) => sum_vector_4_18_port, a(17) => 
                           sum_vector_4_17_port, a(16) => sum_vector_4_16_port,
                           a(15) => sum_vector_4_15_port, a(14) => 
                           sum_vector_4_14_port, a(13) => sum_vector_4_13_port,
                           a(12) => sum_vector_4_12_port, a(11) => 
                           sum_vector_4_11_port, a(10) => sum_vector_4_10_port,
                           a(9) => sum_vector_4_9_port, a(8) => 
                           sum_vector_4_8_port, a(7) => sum_vector_4_7_port, 
                           a(6) => sum_vector_4_6_port, a(5) => 
                           sum_vector_4_5_port, a(4) => sum_vector_4_4_port, 
                           a(3) => sum_vector_4_3_port, a(2) => 
                           sum_vector_4_2_port, a(1) => sum_vector_4_1_port, 
                           a(0) => sum_vector_4_0_port, b(31) => 
                           sum_vector_5_31_port, b(30) => sum_vector_5_30_port,
                           b(29) => sum_vector_5_29_port, b(28) => 
                           sum_vector_5_28_port, b(27) => sum_vector_5_27_port,
                           b(26) => sum_vector_5_26_port, b(25) => 
                           sum_vector_5_25_port, b(24) => sum_vector_5_24_port,
                           b(23) => sum_vector_5_23_port, b(22) => 
                           sum_vector_5_22_port, b(21) => sum_vector_5_21_port,
                           b(20) => sum_vector_5_20_port, b(19) => 
                           sum_vector_5_19_port, b(18) => sum_vector_5_18_port,
                           b(17) => sum_vector_5_17_port, b(16) => 
                           sum_vector_5_16_port, b(15) => sum_vector_5_15_port,
                           b(14) => sum_vector_5_14_port, b(13) => 
                           sum_vector_5_13_port, b(12) => sum_vector_5_12_port,
                           b(11) => sum_vector_5_11_port, b(10) => 
                           sum_vector_5_10_port, b(9) => sum_vector_5_9_port, 
                           b(8) => sum_vector_5_8_port, b(7) => 
                           sum_vector_5_7_port, b(6) => sum_vector_5_6_port, 
                           b(5) => sum_vector_5_5_port, b(4) => 
                           sum_vector_5_4_port, b(3) => sum_vector_5_3_port, 
                           b(2) => sum_vector_5_2_port, b(1) => 
                           sum_vector_5_1_port, b(0) => sum_vector_5_0_port, c 
                           => n_1222, s(31) => sum_vector_6_31_port, s(30) => 
                           sum_vector_6_30_port, s(29) => sum_vector_6_29_port,
                           s(28) => sum_vector_6_28_port, s(27) => 
                           sum_vector_6_27_port, s(26) => sum_vector_6_26_port,
                           s(25) => sum_vector_6_25_port, s(24) => 
                           sum_vector_6_24_port, s(23) => sum_vector_6_23_port,
                           s(22) => sum_vector_6_22_port, s(21) => 
                           sum_vector_6_21_port, s(20) => sum_vector_6_20_port,
                           s(19) => sum_vector_6_19_port, s(18) => 
                           sum_vector_6_18_port, s(17) => sum_vector_6_17_port,
                           s(16) => sum_vector_6_16_port, s(15) => 
                           sum_vector_6_15_port, s(14) => sum_vector_6_14_port,
                           s(13) => sum_vector_6_13_port, s(12) => 
                           sum_vector_6_12_port, s(11) => sum_vector_6_11_port,
                           s(10) => sum_vector_6_10_port, s(9) => 
                           sum_vector_6_9_port, s(8) => sum_vector_6_8_port, 
                           s(7) => sum_vector_6_7_port, s(6) => 
                           sum_vector_6_6_port, s(5) => sum_vector_6_5_port, 
                           s(4) => sum_vector_6_4_port, s(3) => 
                           sum_vector_6_3_port, s(2) => sum_vector_6_2_port, 
                           s(1) => sum_vector_6_1_port, s(0) => 
                           sum_vector_6_0_port);
   shn_4 : shift_NBIT32_SHIFT4 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_4_31_port, pos_a(30) => 
                           pos_av_4_30_port, pos_a(29) => pos_av_4_29_port, 
                           pos_a(28) => pos_av_4_28_port, pos_a(27) => 
                           pos_av_4_27_port, pos_a(26) => pos_av_4_26_port, 
                           pos_a(25) => pos_av_4_25_port, pos_a(24) => 
                           pos_av_4_24_port, pos_a(23) => pos_av_4_23_port, 
                           pos_a(22) => pos_av_4_22_port, pos_a(21) => 
                           pos_av_4_21_port, pos_a(20) => pos_av_4_20_port, 
                           pos_a(19) => pos_av_4_19_port, pos_a(18) => 
                           pos_av_4_18_port, pos_a(17) => pos_av_4_17_port, 
                           pos_a(16) => pos_av_4_16_port, pos_a(15) => 
                           pos_av_4_15_port, pos_a(14) => pos_av_4_14_port, 
                           pos_a(13) => pos_av_4_13_port, pos_a(12) => 
                           pos_av_4_12_port, pos_a(11) => pos_av_4_11_port, 
                           pos_a(10) => pos_av_4_10_port, pos_a(9) => 
                           pos_av_4_9_port, pos_a(8) => pos_av_4_8_port, 
                           pos_a(7) => n_1223, pos_a(6) => n_1224, pos_a(5) => 
                           n_1225, pos_a(4) => n_1226, pos_a(3) => n_1227, 
                           pos_a(2) => n_1228, pos_a(1) => n_1229, pos_a(0) => 
                           n_1230, neg_a(31) => neg_av_4_31_port, neg_a(30) => 
                           neg_av_4_30_port, neg_a(29) => neg_av_4_29_port, 
                           neg_a(28) => neg_av_4_28_port, neg_a(27) => 
                           neg_av_4_27_port, neg_a(26) => neg_av_4_26_port, 
                           neg_a(25) => neg_av_4_25_port, neg_a(24) => 
                           neg_av_4_24_port, neg_a(23) => neg_av_4_23_port, 
                           neg_a(22) => neg_av_4_22_port, neg_a(21) => 
                           neg_av_4_21_port, neg_a(20) => neg_av_4_20_port, 
                           neg_a(19) => neg_av_4_19_port, neg_a(18) => 
                           neg_av_4_18_port, neg_a(17) => neg_av_4_17_port, 
                           neg_a(16) => neg_av_4_16_port, neg_a(15) => 
                           neg_av_4_15_port, neg_a(14) => neg_av_4_14_port, 
                           neg_a(13) => neg_av_4_13_port, neg_a(12) => 
                           neg_av_4_12_port, neg_a(11) => neg_av_4_11_port, 
                           neg_a(10) => neg_av_4_10_port, neg_a(9) => 
                           neg_av_4_9_port, neg_a(8) => neg_av_4_8_port, 
                           neg_a(7) => n_1231, neg_a(6) => n_1232, neg_a(5) => 
                           n_1233, neg_a(4) => n_1234, neg_a(3) => n_1235, 
                           neg_a(2) => n_1236, neg_a(1) => n_1237, neg_a(0) => 
                           n_1238, pos_2a(31) => pos_2av_4_31_port, pos_2a(30) 
                           => pos_2av_4_30_port, pos_2a(29) => 
                           pos_2av_4_29_port, pos_2a(28) => pos_2av_4_28_port, 
                           pos_2a(27) => pos_2av_4_27_port, pos_2a(26) => 
                           pos_2av_4_26_port, pos_2a(25) => pos_2av_4_25_port, 
                           pos_2a(24) => pos_2av_4_24_port, pos_2a(23) => 
                           pos_2av_4_23_port, pos_2a(22) => pos_2av_4_22_port, 
                           pos_2a(21) => pos_2av_4_21_port, pos_2a(20) => 
                           pos_2av_4_20_port, pos_2a(19) => pos_2av_4_19_port, 
                           pos_2a(18) => pos_2av_4_18_port, pos_2a(17) => 
                           pos_2av_4_17_port, pos_2a(16) => pos_2av_4_16_port, 
                           pos_2a(15) => pos_2av_4_15_port, pos_2a(14) => 
                           pos_2av_4_14_port, pos_2a(13) => pos_2av_4_13_port, 
                           pos_2a(12) => pos_2av_4_12_port, pos_2a(11) => 
                           pos_2av_4_11_port, pos_2a(10) => pos_2av_4_10_port, 
                           pos_2a(9) => pos_2av_4_9_port, pos_2a(8) => n_1239, 
                           pos_2a(7) => n_1240, pos_2a(6) => n_1241, pos_2a(5) 
                           => n_1242, pos_2a(4) => n_1243, pos_2a(3) => n_1244,
                           pos_2a(2) => n_1245, pos_2a(1) => n_1246, pos_2a(0) 
                           => n_1247, neg_2a(31) => neg_2av_4_31_port, 
                           neg_2a(30) => neg_2av_4_30_port, neg_2a(29) => 
                           neg_2av_4_29_port, neg_2a(28) => neg_2av_4_28_port, 
                           neg_2a(27) => neg_2av_4_27_port, neg_2a(26) => 
                           neg_2av_4_26_port, neg_2a(25) => neg_2av_4_25_port, 
                           neg_2a(24) => neg_2av_4_24_port, neg_2a(23) => 
                           neg_2av_4_23_port, neg_2a(22) => neg_2av_4_22_port, 
                           neg_2a(21) => neg_2av_4_21_port, neg_2a(20) => 
                           neg_2av_4_20_port, neg_2a(19) => neg_2av_4_19_port, 
                           neg_2a(18) => neg_2av_4_18_port, neg_2a(17) => 
                           neg_2av_4_17_port, neg_2a(16) => neg_2av_4_16_port, 
                           neg_2a(15) => neg_2av_4_15_port, neg_2a(14) => 
                           neg_2av_4_14_port, neg_2a(13) => neg_2av_4_13_port, 
                           neg_2a(12) => neg_2av_4_12_port, neg_2a(11) => 
                           neg_2av_4_11_port, neg_2a(10) => neg_2av_4_10_port, 
                           neg_2a(9) => neg_2av_4_9_port, neg_2a(8) => n_1248, 
                           neg_2a(7) => n_1249, neg_2a(6) => n_1250, neg_2a(5) 
                           => n_1251, neg_2a(4) => n_1252, neg_2a(3) => n_1253,
                           neg_2a(2) => n_1254, neg_2a(1) => n_1255, neg_2a(0) 
                           => n_1256);
   vpn_4 : vp_NBIT32_4 port map( pos_a(31) => pos_av_4_31_port, pos_a(30) => 
                           pos_av_4_30_port, pos_a(29) => pos_av_4_29_port, 
                           pos_a(28) => pos_av_4_28_port, pos_a(27) => 
                           pos_av_4_27_port, pos_a(26) => pos_av_4_26_port, 
                           pos_a(25) => pos_av_4_25_port, pos_a(24) => 
                           pos_av_4_24_port, pos_a(23) => pos_av_4_23_port, 
                           pos_a(22) => pos_av_4_22_port, pos_a(21) => 
                           pos_av_4_21_port, pos_a(20) => pos_av_4_20_port, 
                           pos_a(19) => pos_av_4_19_port, pos_a(18) => 
                           pos_av_4_18_port, pos_a(17) => pos_av_4_17_port, 
                           pos_a(16) => pos_av_4_16_port, pos_a(15) => 
                           pos_av_4_15_port, pos_a(14) => pos_av_4_14_port, 
                           pos_a(13) => pos_av_4_13_port, pos_a(12) => 
                           pos_av_4_12_port, pos_a(11) => pos_av_4_11_port, 
                           pos_a(10) => pos_av_4_10_port, pos_a(9) => 
                           pos_av_4_9_port, pos_a(8) => pos_av_4_8_port, 
                           pos_a(7) => pos_av_4_7_port, pos_a(6) => 
                           pos_av_4_6_port, pos_a(5) => pos_av_4_5_port, 
                           pos_a(4) => pos_av_4_4_port, pos_a(3) => 
                           pos_av_4_3_port, pos_a(2) => pos_av_4_2_port, 
                           pos_a(1) => pos_av_4_1_port, pos_a(0) => 
                           pos_av_4_0_port, neg_a(31) => neg_av_4_31_port, 
                           neg_a(30) => neg_av_4_30_port, neg_a(29) => 
                           neg_av_4_29_port, neg_a(28) => neg_av_4_28_port, 
                           neg_a(27) => neg_av_4_27_port, neg_a(26) => 
                           neg_av_4_26_port, neg_a(25) => neg_av_4_25_port, 
                           neg_a(24) => neg_av_4_24_port, neg_a(23) => 
                           neg_av_4_23_port, neg_a(22) => neg_av_4_22_port, 
                           neg_a(21) => neg_av_4_21_port, neg_a(20) => 
                           neg_av_4_20_port, neg_a(19) => neg_av_4_19_port, 
                           neg_a(18) => neg_av_4_18_port, neg_a(17) => 
                           neg_av_4_17_port, neg_a(16) => neg_av_4_16_port, 
                           neg_a(15) => neg_av_4_15_port, neg_a(14) => 
                           neg_av_4_14_port, neg_a(13) => neg_av_4_13_port, 
                           neg_a(12) => neg_av_4_12_port, neg_a(11) => 
                           neg_av_4_11_port, neg_a(10) => neg_av_4_10_port, 
                           neg_a(9) => neg_av_4_9_port, neg_a(8) => 
                           neg_av_4_8_port, neg_a(7) => neg_av_4_7_port, 
                           neg_a(6) => neg_av_4_6_port, neg_a(5) => 
                           neg_av_4_5_port, neg_a(4) => neg_av_4_4_port, 
                           neg_a(3) => neg_av_4_3_port, neg_a(2) => 
                           neg_av_4_2_port, neg_a(1) => neg_av_4_1_port, 
                           neg_a(0) => neg_av_4_0_port, pos_2a(31) => 
                           pos_2av_4_31_port, pos_2a(30) => pos_2av_4_30_port, 
                           pos_2a(29) => pos_2av_4_29_port, pos_2a(28) => 
                           pos_2av_4_28_port, pos_2a(27) => pos_2av_4_27_port, 
                           pos_2a(26) => pos_2av_4_26_port, pos_2a(25) => 
                           pos_2av_4_25_port, pos_2a(24) => pos_2av_4_24_port, 
                           pos_2a(23) => pos_2av_4_23_port, pos_2a(22) => 
                           pos_2av_4_22_port, pos_2a(21) => pos_2av_4_21_port, 
                           pos_2a(20) => pos_2av_4_20_port, pos_2a(19) => 
                           pos_2av_4_19_port, pos_2a(18) => pos_2av_4_18_port, 
                           pos_2a(17) => pos_2av_4_17_port, pos_2a(16) => 
                           pos_2av_4_16_port, pos_2a(15) => pos_2av_4_15_port, 
                           pos_2a(14) => pos_2av_4_14_port, pos_2a(13) => 
                           pos_2av_4_13_port, pos_2a(12) => pos_2av_4_12_port, 
                           pos_2a(11) => pos_2av_4_11_port, pos_2a(10) => 
                           pos_2av_4_10_port, pos_2a(9) => pos_2av_4_9_port, 
                           pos_2a(8) => pos_2av_4_8_port, pos_2a(7) => 
                           pos_2av_4_7_port, pos_2a(6) => pos_2av_4_6_port, 
                           pos_2a(5) => pos_2av_4_5_port, pos_2a(4) => 
                           pos_2av_4_4_port, pos_2a(3) => pos_2av_4_3_port, 
                           pos_2a(2) => pos_2av_4_2_port, pos_2a(1) => 
                           pos_2av_4_1_port, pos_2a(0) => pos_2av_4_0_port, 
                           neg_2a(31) => neg_2av_4_31_port, neg_2a(30) => 
                           neg_2av_4_30_port, neg_2a(29) => neg_2av_4_29_port, 
                           neg_2a(28) => neg_2av_4_28_port, neg_2a(27) => 
                           neg_2av_4_27_port, neg_2a(26) => neg_2av_4_26_port, 
                           neg_2a(25) => neg_2av_4_25_port, neg_2a(24) => 
                           neg_2av_4_24_port, neg_2a(23) => neg_2av_4_23_port, 
                           neg_2a(22) => neg_2av_4_22_port, neg_2a(21) => 
                           neg_2av_4_21_port, neg_2a(20) => neg_2av_4_20_port, 
                           neg_2a(19) => neg_2av_4_19_port, neg_2a(18) => 
                           neg_2av_4_18_port, neg_2a(17) => neg_2av_4_17_port, 
                           neg_2a(16) => neg_2av_4_16_port, neg_2a(15) => 
                           neg_2av_4_15_port, neg_2a(14) => neg_2av_4_14_port, 
                           neg_2a(13) => neg_2av_4_13_port, neg_2a(12) => 
                           neg_2av_4_12_port, neg_2a(11) => neg_2av_4_11_port, 
                           neg_2a(10) => neg_2av_4_10_port, neg_2a(9) => 
                           neg_2av_4_9_port, neg_2a(8) => neg_2av_4_8_port, 
                           neg_2a(7) => neg_2av_4_7_port, neg_2a(6) => 
                           neg_2av_4_6_port, neg_2a(5) => neg_2av_4_5_port, 
                           neg_2a(4) => neg_2av_4_4_port, neg_2a(3) => 
                           neg_2av_4_3_port, neg_2a(2) => neg_2av_4_2_port, 
                           neg_2a(1) => neg_2av_4_1_port, neg_2a(0) => 
                           neg_2av_4_0_port, sel(2) => b(9), sel(1) => b(8), 
                           sel(0) => b(7), s_out(31) => sum_vector_7_31_port, 
                           s_out(30) => sum_vector_7_30_port, s_out(29) => 
                           sum_vector_7_29_port, s_out(28) => 
                           sum_vector_7_28_port, s_out(27) => 
                           sum_vector_7_27_port, s_out(26) => 
                           sum_vector_7_26_port, s_out(25) => 
                           sum_vector_7_25_port, s_out(24) => 
                           sum_vector_7_24_port, s_out(23) => 
                           sum_vector_7_23_port, s_out(22) => 
                           sum_vector_7_22_port, s_out(21) => 
                           sum_vector_7_21_port, s_out(20) => 
                           sum_vector_7_20_port, s_out(19) => 
                           sum_vector_7_19_port, s_out(18) => 
                           sum_vector_7_18_port, s_out(17) => 
                           sum_vector_7_17_port, s_out(16) => 
                           sum_vector_7_16_port, s_out(15) => 
                           sum_vector_7_15_port, s_out(14) => 
                           sum_vector_7_14_port, s_out(13) => 
                           sum_vector_7_13_port, s_out(12) => 
                           sum_vector_7_12_port, s_out(11) => 
                           sum_vector_7_11_port, s_out(10) => 
                           sum_vector_7_10_port, s_out(9) => 
                           sum_vector_7_9_port, s_out(8) => sum_vector_7_8_port
                           , s_out(7) => sum_vector_7_7_port, s_out(6) => 
                           sum_vector_7_6_port, s_out(5) => sum_vector_7_5_port
                           , s_out(4) => sum_vector_7_4_port, s_out(3) => 
                           sum_vector_7_3_port, s_out(2) => sum_vector_7_2_port
                           , s_out(1) => sum_vector_7_1_port, s_out(0) => 
                           sum_vector_7_0_port);
   sumn_4 : rca_signed_NBIT32_4 port map( a(31) => sum_vector_6_31_port, a(30) 
                           => sum_vector_6_30_port, a(29) => 
                           sum_vector_6_29_port, a(28) => sum_vector_6_28_port,
                           a(27) => sum_vector_6_27_port, a(26) => 
                           sum_vector_6_26_port, a(25) => sum_vector_6_25_port,
                           a(24) => sum_vector_6_24_port, a(23) => 
                           sum_vector_6_23_port, a(22) => sum_vector_6_22_port,
                           a(21) => sum_vector_6_21_port, a(20) => 
                           sum_vector_6_20_port, a(19) => sum_vector_6_19_port,
                           a(18) => sum_vector_6_18_port, a(17) => 
                           sum_vector_6_17_port, a(16) => sum_vector_6_16_port,
                           a(15) => sum_vector_6_15_port, a(14) => 
                           sum_vector_6_14_port, a(13) => sum_vector_6_13_port,
                           a(12) => sum_vector_6_12_port, a(11) => 
                           sum_vector_6_11_port, a(10) => sum_vector_6_10_port,
                           a(9) => sum_vector_6_9_port, a(8) => 
                           sum_vector_6_8_port, a(7) => sum_vector_6_7_port, 
                           a(6) => sum_vector_6_6_port, a(5) => 
                           sum_vector_6_5_port, a(4) => sum_vector_6_4_port, 
                           a(3) => sum_vector_6_3_port, a(2) => 
                           sum_vector_6_2_port, a(1) => sum_vector_6_1_port, 
                           a(0) => sum_vector_6_0_port, b(31) => 
                           sum_vector_7_31_port, b(30) => sum_vector_7_30_port,
                           b(29) => sum_vector_7_29_port, b(28) => 
                           sum_vector_7_28_port, b(27) => sum_vector_7_27_port,
                           b(26) => sum_vector_7_26_port, b(25) => 
                           sum_vector_7_25_port, b(24) => sum_vector_7_24_port,
                           b(23) => sum_vector_7_23_port, b(22) => 
                           sum_vector_7_22_port, b(21) => sum_vector_7_21_port,
                           b(20) => sum_vector_7_20_port, b(19) => 
                           sum_vector_7_19_port, b(18) => sum_vector_7_18_port,
                           b(17) => sum_vector_7_17_port, b(16) => 
                           sum_vector_7_16_port, b(15) => sum_vector_7_15_port,
                           b(14) => sum_vector_7_14_port, b(13) => 
                           sum_vector_7_13_port, b(12) => sum_vector_7_12_port,
                           b(11) => sum_vector_7_11_port, b(10) => 
                           sum_vector_7_10_port, b(9) => sum_vector_7_9_port, 
                           b(8) => sum_vector_7_8_port, b(7) => 
                           sum_vector_7_7_port, b(6) => sum_vector_7_6_port, 
                           b(5) => sum_vector_7_5_port, b(4) => 
                           sum_vector_7_4_port, b(3) => sum_vector_7_3_port, 
                           b(2) => sum_vector_7_2_port, b(1) => 
                           sum_vector_7_1_port, b(0) => sum_vector_7_0_port, c 
                           => n_1257, s(31) => sum_vector_8_31_port, s(30) => 
                           sum_vector_8_30_port, s(29) => sum_vector_8_29_port,
                           s(28) => sum_vector_8_28_port, s(27) => 
                           sum_vector_8_27_port, s(26) => sum_vector_8_26_port,
                           s(25) => sum_vector_8_25_port, s(24) => 
                           sum_vector_8_24_port, s(23) => sum_vector_8_23_port,
                           s(22) => sum_vector_8_22_port, s(21) => 
                           sum_vector_8_21_port, s(20) => sum_vector_8_20_port,
                           s(19) => sum_vector_8_19_port, s(18) => 
                           sum_vector_8_18_port, s(17) => sum_vector_8_17_port,
                           s(16) => sum_vector_8_16_port, s(15) => 
                           sum_vector_8_15_port, s(14) => sum_vector_8_14_port,
                           s(13) => sum_vector_8_13_port, s(12) => 
                           sum_vector_8_12_port, s(11) => sum_vector_8_11_port,
                           s(10) => sum_vector_8_10_port, s(9) => 
                           sum_vector_8_9_port, s(8) => sum_vector_8_8_port, 
                           s(7) => sum_vector_8_7_port, s(6) => 
                           sum_vector_8_6_port, s(5) => sum_vector_8_5_port, 
                           s(4) => sum_vector_8_4_port, s(3) => 
                           sum_vector_8_3_port, s(2) => sum_vector_8_2_port, 
                           s(1) => sum_vector_8_1_port, s(0) => 
                           sum_vector_8_0_port);
   shn_5 : shift_NBIT32_SHIFT5 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_5_31_port, pos_a(30) => 
                           pos_av_5_30_port, pos_a(29) => pos_av_5_29_port, 
                           pos_a(28) => pos_av_5_28_port, pos_a(27) => 
                           pos_av_5_27_port, pos_a(26) => pos_av_5_26_port, 
                           pos_a(25) => pos_av_5_25_port, pos_a(24) => 
                           pos_av_5_24_port, pos_a(23) => pos_av_5_23_port, 
                           pos_a(22) => pos_av_5_22_port, pos_a(21) => 
                           pos_av_5_21_port, pos_a(20) => pos_av_5_20_port, 
                           pos_a(19) => pos_av_5_19_port, pos_a(18) => 
                           pos_av_5_18_port, pos_a(17) => pos_av_5_17_port, 
                           pos_a(16) => pos_av_5_16_port, pos_a(15) => 
                           pos_av_5_15_port, pos_a(14) => pos_av_5_14_port, 
                           pos_a(13) => pos_av_5_13_port, pos_a(12) => 
                           pos_av_5_12_port, pos_a(11) => pos_av_5_11_port, 
                           pos_a(10) => pos_av_5_10_port, pos_a(9) => n_1258, 
                           pos_a(8) => n_1259, pos_a(7) => n_1260, pos_a(6) => 
                           n_1261, pos_a(5) => n_1262, pos_a(4) => n_1263, 
                           pos_a(3) => n_1264, pos_a(2) => n_1265, pos_a(1) => 
                           n_1266, pos_a(0) => n_1267, neg_a(31) => 
                           neg_av_5_31_port, neg_a(30) => neg_av_5_30_port, 
                           neg_a(29) => neg_av_5_29_port, neg_a(28) => 
                           neg_av_5_28_port, neg_a(27) => neg_av_5_27_port, 
                           neg_a(26) => neg_av_5_26_port, neg_a(25) => 
                           neg_av_5_25_port, neg_a(24) => neg_av_5_24_port, 
                           neg_a(23) => neg_av_5_23_port, neg_a(22) => 
                           neg_av_5_22_port, neg_a(21) => neg_av_5_21_port, 
                           neg_a(20) => neg_av_5_20_port, neg_a(19) => 
                           neg_av_5_19_port, neg_a(18) => neg_av_5_18_port, 
                           neg_a(17) => neg_av_5_17_port, neg_a(16) => 
                           neg_av_5_16_port, neg_a(15) => neg_av_5_15_port, 
                           neg_a(14) => neg_av_5_14_port, neg_a(13) => 
                           neg_av_5_13_port, neg_a(12) => neg_av_5_12_port, 
                           neg_a(11) => neg_av_5_11_port, neg_a(10) => 
                           neg_av_5_10_port, neg_a(9) => n_1268, neg_a(8) => 
                           n_1269, neg_a(7) => n_1270, neg_a(6) => n_1271, 
                           neg_a(5) => n_1272, neg_a(4) => n_1273, neg_a(3) => 
                           n_1274, neg_a(2) => n_1275, neg_a(1) => n_1276, 
                           neg_a(0) => n_1277, pos_2a(31) => pos_2av_5_31_port,
                           pos_2a(30) => pos_2av_5_30_port, pos_2a(29) => 
                           pos_2av_5_29_port, pos_2a(28) => pos_2av_5_28_port, 
                           pos_2a(27) => pos_2av_5_27_port, pos_2a(26) => 
                           pos_2av_5_26_port, pos_2a(25) => pos_2av_5_25_port, 
                           pos_2a(24) => pos_2av_5_24_port, pos_2a(23) => 
                           pos_2av_5_23_port, pos_2a(22) => pos_2av_5_22_port, 
                           pos_2a(21) => pos_2av_5_21_port, pos_2a(20) => 
                           pos_2av_5_20_port, pos_2a(19) => pos_2av_5_19_port, 
                           pos_2a(18) => pos_2av_5_18_port, pos_2a(17) => 
                           pos_2av_5_17_port, pos_2a(16) => pos_2av_5_16_port, 
                           pos_2a(15) => pos_2av_5_15_port, pos_2a(14) => 
                           pos_2av_5_14_port, pos_2a(13) => pos_2av_5_13_port, 
                           pos_2a(12) => pos_2av_5_12_port, pos_2a(11) => 
                           pos_2av_5_11_port, pos_2a(10) => n_1278, pos_2a(9) 
                           => n_1279, pos_2a(8) => n_1280, pos_2a(7) => n_1281,
                           pos_2a(6) => n_1282, pos_2a(5) => n_1283, pos_2a(4) 
                           => n_1284, pos_2a(3) => n_1285, pos_2a(2) => n_1286,
                           pos_2a(1) => n_1287, pos_2a(0) => n_1288, neg_2a(31)
                           => neg_2av_5_31_port, neg_2a(30) => 
                           neg_2av_5_30_port, neg_2a(29) => neg_2av_5_29_port, 
                           neg_2a(28) => neg_2av_5_28_port, neg_2a(27) => 
                           neg_2av_5_27_port, neg_2a(26) => neg_2av_5_26_port, 
                           neg_2a(25) => neg_2av_5_25_port, neg_2a(24) => 
                           neg_2av_5_24_port, neg_2a(23) => neg_2av_5_23_port, 
                           neg_2a(22) => neg_2av_5_22_port, neg_2a(21) => 
                           neg_2av_5_21_port, neg_2a(20) => neg_2av_5_20_port, 
                           neg_2a(19) => neg_2av_5_19_port, neg_2a(18) => 
                           neg_2av_5_18_port, neg_2a(17) => neg_2av_5_17_port, 
                           neg_2a(16) => neg_2av_5_16_port, neg_2a(15) => 
                           neg_2av_5_15_port, neg_2a(14) => neg_2av_5_14_port, 
                           neg_2a(13) => neg_2av_5_13_port, neg_2a(12) => 
                           neg_2av_5_12_port, neg_2a(11) => neg_2av_5_11_port, 
                           neg_2a(10) => n_1289, neg_2a(9) => n_1290, neg_2a(8)
                           => n_1291, neg_2a(7) => n_1292, neg_2a(6) => n_1293,
                           neg_2a(5) => n_1294, neg_2a(4) => n_1295, neg_2a(3) 
                           => n_1296, neg_2a(2) => n_1297, neg_2a(1) => n_1298,
                           neg_2a(0) => n_1299);
   vpn_5 : vp_NBIT32_3 port map( pos_a(31) => pos_av_5_31_port, pos_a(30) => 
                           pos_av_5_30_port, pos_a(29) => pos_av_5_29_port, 
                           pos_a(28) => pos_av_5_28_port, pos_a(27) => 
                           pos_av_5_27_port, pos_a(26) => pos_av_5_26_port, 
                           pos_a(25) => pos_av_5_25_port, pos_a(24) => 
                           pos_av_5_24_port, pos_a(23) => pos_av_5_23_port, 
                           pos_a(22) => pos_av_5_22_port, pos_a(21) => 
                           pos_av_5_21_port, pos_a(20) => pos_av_5_20_port, 
                           pos_a(19) => pos_av_5_19_port, pos_a(18) => 
                           pos_av_5_18_port, pos_a(17) => pos_av_5_17_port, 
                           pos_a(16) => pos_av_5_16_port, pos_a(15) => 
                           pos_av_5_15_port, pos_a(14) => pos_av_5_14_port, 
                           pos_a(13) => pos_av_5_13_port, pos_a(12) => 
                           pos_av_5_12_port, pos_a(11) => pos_av_5_11_port, 
                           pos_a(10) => pos_av_5_10_port, pos_a(9) => 
                           pos_av_5_9_port, pos_a(8) => pos_av_5_8_port, 
                           pos_a(7) => pos_av_5_7_port, pos_a(6) => 
                           pos_av_5_6_port, pos_a(5) => pos_av_5_5_port, 
                           pos_a(4) => pos_av_5_4_port, pos_a(3) => 
                           pos_av_5_3_port, pos_a(2) => pos_av_5_2_port, 
                           pos_a(1) => pos_av_5_1_port, pos_a(0) => 
                           pos_av_5_0_port, neg_a(31) => neg_av_5_31_port, 
                           neg_a(30) => neg_av_5_30_port, neg_a(29) => 
                           neg_av_5_29_port, neg_a(28) => neg_av_5_28_port, 
                           neg_a(27) => neg_av_5_27_port, neg_a(26) => 
                           neg_av_5_26_port, neg_a(25) => neg_av_5_25_port, 
                           neg_a(24) => neg_av_5_24_port, neg_a(23) => 
                           neg_av_5_23_port, neg_a(22) => neg_av_5_22_port, 
                           neg_a(21) => neg_av_5_21_port, neg_a(20) => 
                           neg_av_5_20_port, neg_a(19) => neg_av_5_19_port, 
                           neg_a(18) => neg_av_5_18_port, neg_a(17) => 
                           neg_av_5_17_port, neg_a(16) => neg_av_5_16_port, 
                           neg_a(15) => neg_av_5_15_port, neg_a(14) => 
                           neg_av_5_14_port, neg_a(13) => neg_av_5_13_port, 
                           neg_a(12) => neg_av_5_12_port, neg_a(11) => 
                           neg_av_5_11_port, neg_a(10) => neg_av_5_10_port, 
                           neg_a(9) => neg_av_5_9_port, neg_a(8) => 
                           neg_av_5_8_port, neg_a(7) => neg_av_5_7_port, 
                           neg_a(6) => neg_av_5_6_port, neg_a(5) => 
                           neg_av_5_5_port, neg_a(4) => neg_av_5_4_port, 
                           neg_a(3) => neg_av_5_3_port, neg_a(2) => 
                           neg_av_5_2_port, neg_a(1) => neg_av_5_1_port, 
                           neg_a(0) => neg_av_5_0_port, pos_2a(31) => 
                           pos_2av_5_31_port, pos_2a(30) => pos_2av_5_30_port, 
                           pos_2a(29) => pos_2av_5_29_port, pos_2a(28) => 
                           pos_2av_5_28_port, pos_2a(27) => pos_2av_5_27_port, 
                           pos_2a(26) => pos_2av_5_26_port, pos_2a(25) => 
                           pos_2av_5_25_port, pos_2a(24) => pos_2av_5_24_port, 
                           pos_2a(23) => pos_2av_5_23_port, pos_2a(22) => 
                           pos_2av_5_22_port, pos_2a(21) => pos_2av_5_21_port, 
                           pos_2a(20) => pos_2av_5_20_port, pos_2a(19) => 
                           pos_2av_5_19_port, pos_2a(18) => pos_2av_5_18_port, 
                           pos_2a(17) => pos_2av_5_17_port, pos_2a(16) => 
                           pos_2av_5_16_port, pos_2a(15) => pos_2av_5_15_port, 
                           pos_2a(14) => pos_2av_5_14_port, pos_2a(13) => 
                           pos_2av_5_13_port, pos_2a(12) => pos_2av_5_12_port, 
                           pos_2a(11) => pos_2av_5_11_port, pos_2a(10) => 
                           pos_2av_5_10_port, pos_2a(9) => pos_2av_5_9_port, 
                           pos_2a(8) => pos_2av_5_8_port, pos_2a(7) => 
                           pos_2av_5_7_port, pos_2a(6) => pos_2av_5_6_port, 
                           pos_2a(5) => pos_2av_5_5_port, pos_2a(4) => 
                           pos_2av_5_4_port, pos_2a(3) => pos_2av_5_3_port, 
                           pos_2a(2) => pos_2av_5_2_port, pos_2a(1) => 
                           pos_2av_5_1_port, pos_2a(0) => pos_2av_5_0_port, 
                           neg_2a(31) => neg_2av_5_31_port, neg_2a(30) => 
                           neg_2av_5_30_port, neg_2a(29) => neg_2av_5_29_port, 
                           neg_2a(28) => neg_2av_5_28_port, neg_2a(27) => 
                           neg_2av_5_27_port, neg_2a(26) => neg_2av_5_26_port, 
                           neg_2a(25) => neg_2av_5_25_port, neg_2a(24) => 
                           neg_2av_5_24_port, neg_2a(23) => neg_2av_5_23_port, 
                           neg_2a(22) => neg_2av_5_22_port, neg_2a(21) => 
                           neg_2av_5_21_port, neg_2a(20) => neg_2av_5_20_port, 
                           neg_2a(19) => neg_2av_5_19_port, neg_2a(18) => 
                           neg_2av_5_18_port, neg_2a(17) => neg_2av_5_17_port, 
                           neg_2a(16) => neg_2av_5_16_port, neg_2a(15) => 
                           neg_2av_5_15_port, neg_2a(14) => neg_2av_5_14_port, 
                           neg_2a(13) => neg_2av_5_13_port, neg_2a(12) => 
                           neg_2av_5_12_port, neg_2a(11) => neg_2av_5_11_port, 
                           neg_2a(10) => neg_2av_5_10_port, neg_2a(9) => 
                           neg_2av_5_9_port, neg_2a(8) => neg_2av_5_8_port, 
                           neg_2a(7) => neg_2av_5_7_port, neg_2a(6) => 
                           neg_2av_5_6_port, neg_2a(5) => neg_2av_5_5_port, 
                           neg_2a(4) => neg_2av_5_4_port, neg_2a(3) => 
                           neg_2av_5_3_port, neg_2a(2) => neg_2av_5_2_port, 
                           neg_2a(1) => neg_2av_5_1_port, neg_2a(0) => 
                           neg_2av_5_0_port, sel(2) => b(11), sel(1) => b(10), 
                           sel(0) => b(9), s_out(31) => sum_vector_9_31_port, 
                           s_out(30) => sum_vector_9_30_port, s_out(29) => 
                           sum_vector_9_29_port, s_out(28) => 
                           sum_vector_9_28_port, s_out(27) => 
                           sum_vector_9_27_port, s_out(26) => 
                           sum_vector_9_26_port, s_out(25) => 
                           sum_vector_9_25_port, s_out(24) => 
                           sum_vector_9_24_port, s_out(23) => 
                           sum_vector_9_23_port, s_out(22) => 
                           sum_vector_9_22_port, s_out(21) => 
                           sum_vector_9_21_port, s_out(20) => 
                           sum_vector_9_20_port, s_out(19) => 
                           sum_vector_9_19_port, s_out(18) => 
                           sum_vector_9_18_port, s_out(17) => 
                           sum_vector_9_17_port, s_out(16) => 
                           sum_vector_9_16_port, s_out(15) => 
                           sum_vector_9_15_port, s_out(14) => 
                           sum_vector_9_14_port, s_out(13) => 
                           sum_vector_9_13_port, s_out(12) => 
                           sum_vector_9_12_port, s_out(11) => 
                           sum_vector_9_11_port, s_out(10) => 
                           sum_vector_9_10_port, s_out(9) => 
                           sum_vector_9_9_port, s_out(8) => sum_vector_9_8_port
                           , s_out(7) => sum_vector_9_7_port, s_out(6) => 
                           sum_vector_9_6_port, s_out(5) => sum_vector_9_5_port
                           , s_out(4) => sum_vector_9_4_port, s_out(3) => 
                           sum_vector_9_3_port, s_out(2) => sum_vector_9_2_port
                           , s_out(1) => sum_vector_9_1_port, s_out(0) => 
                           sum_vector_9_0_port);
   sumn_5 : rca_signed_NBIT32_3 port map( a(31) => sum_vector_8_31_port, a(30) 
                           => sum_vector_8_30_port, a(29) => 
                           sum_vector_8_29_port, a(28) => sum_vector_8_28_port,
                           a(27) => sum_vector_8_27_port, a(26) => 
                           sum_vector_8_26_port, a(25) => sum_vector_8_25_port,
                           a(24) => sum_vector_8_24_port, a(23) => 
                           sum_vector_8_23_port, a(22) => sum_vector_8_22_port,
                           a(21) => sum_vector_8_21_port, a(20) => 
                           sum_vector_8_20_port, a(19) => sum_vector_8_19_port,
                           a(18) => sum_vector_8_18_port, a(17) => 
                           sum_vector_8_17_port, a(16) => sum_vector_8_16_port,
                           a(15) => sum_vector_8_15_port, a(14) => 
                           sum_vector_8_14_port, a(13) => sum_vector_8_13_port,
                           a(12) => sum_vector_8_12_port, a(11) => 
                           sum_vector_8_11_port, a(10) => sum_vector_8_10_port,
                           a(9) => sum_vector_8_9_port, a(8) => 
                           sum_vector_8_8_port, a(7) => sum_vector_8_7_port, 
                           a(6) => sum_vector_8_6_port, a(5) => 
                           sum_vector_8_5_port, a(4) => sum_vector_8_4_port, 
                           a(3) => sum_vector_8_3_port, a(2) => 
                           sum_vector_8_2_port, a(1) => sum_vector_8_1_port, 
                           a(0) => sum_vector_8_0_port, b(31) => 
                           sum_vector_9_31_port, b(30) => sum_vector_9_30_port,
                           b(29) => sum_vector_9_29_port, b(28) => 
                           sum_vector_9_28_port, b(27) => sum_vector_9_27_port,
                           b(26) => sum_vector_9_26_port, b(25) => 
                           sum_vector_9_25_port, b(24) => sum_vector_9_24_port,
                           b(23) => sum_vector_9_23_port, b(22) => 
                           sum_vector_9_22_port, b(21) => sum_vector_9_21_port,
                           b(20) => sum_vector_9_20_port, b(19) => 
                           sum_vector_9_19_port, b(18) => sum_vector_9_18_port,
                           b(17) => sum_vector_9_17_port, b(16) => 
                           sum_vector_9_16_port, b(15) => sum_vector_9_15_port,
                           b(14) => sum_vector_9_14_port, b(13) => 
                           sum_vector_9_13_port, b(12) => sum_vector_9_12_port,
                           b(11) => sum_vector_9_11_port, b(10) => 
                           sum_vector_9_10_port, b(9) => sum_vector_9_9_port, 
                           b(8) => sum_vector_9_8_port, b(7) => 
                           sum_vector_9_7_port, b(6) => sum_vector_9_6_port, 
                           b(5) => sum_vector_9_5_port, b(4) => 
                           sum_vector_9_4_port, b(3) => sum_vector_9_3_port, 
                           b(2) => sum_vector_9_2_port, b(1) => 
                           sum_vector_9_1_port, b(0) => sum_vector_9_0_port, c 
                           => n_1300, s(31) => sum_vector_10_31_port, s(30) => 
                           sum_vector_10_30_port, s(29) => 
                           sum_vector_10_29_port, s(28) => 
                           sum_vector_10_28_port, s(27) => 
                           sum_vector_10_27_port, s(26) => 
                           sum_vector_10_26_port, s(25) => 
                           sum_vector_10_25_port, s(24) => 
                           sum_vector_10_24_port, s(23) => 
                           sum_vector_10_23_port, s(22) => 
                           sum_vector_10_22_port, s(21) => 
                           sum_vector_10_21_port, s(20) => 
                           sum_vector_10_20_port, s(19) => 
                           sum_vector_10_19_port, s(18) => 
                           sum_vector_10_18_port, s(17) => 
                           sum_vector_10_17_port, s(16) => 
                           sum_vector_10_16_port, s(15) => 
                           sum_vector_10_15_port, s(14) => 
                           sum_vector_10_14_port, s(13) => 
                           sum_vector_10_13_port, s(12) => 
                           sum_vector_10_12_port, s(11) => 
                           sum_vector_10_11_port, s(10) => 
                           sum_vector_10_10_port, s(9) => sum_vector_10_9_port,
                           s(8) => sum_vector_10_8_port, s(7) => 
                           sum_vector_10_7_port, s(6) => sum_vector_10_6_port, 
                           s(5) => sum_vector_10_5_port, s(4) => 
                           sum_vector_10_4_port, s(3) => sum_vector_10_3_port, 
                           s(2) => sum_vector_10_2_port, s(1) => 
                           sum_vector_10_1_port, s(0) => sum_vector_10_0_port);
   shn_6 : shift_NBIT32_SHIFT6 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_6_31_port, pos_a(30) => 
                           pos_av_6_30_port, pos_a(29) => pos_av_6_29_port, 
                           pos_a(28) => pos_av_6_28_port, pos_a(27) => 
                           pos_av_6_27_port, pos_a(26) => pos_av_6_26_port, 
                           pos_a(25) => pos_av_6_25_port, pos_a(24) => 
                           pos_av_6_24_port, pos_a(23) => pos_av_6_23_port, 
                           pos_a(22) => pos_av_6_22_port, pos_a(21) => 
                           pos_av_6_21_port, pos_a(20) => pos_av_6_20_port, 
                           pos_a(19) => pos_av_6_19_port, pos_a(18) => 
                           pos_av_6_18_port, pos_a(17) => pos_av_6_17_port, 
                           pos_a(16) => pos_av_6_16_port, pos_a(15) => 
                           pos_av_6_15_port, pos_a(14) => pos_av_6_14_port, 
                           pos_a(13) => pos_av_6_13_port, pos_a(12) => 
                           pos_av_6_12_port, pos_a(11) => n_1301, pos_a(10) => 
                           n_1302, pos_a(9) => n_1303, pos_a(8) => n_1304, 
                           pos_a(7) => n_1305, pos_a(6) => n_1306, pos_a(5) => 
                           n_1307, pos_a(4) => n_1308, pos_a(3) => n_1309, 
                           pos_a(2) => n_1310, pos_a(1) => n_1311, pos_a(0) => 
                           n_1312, neg_a(31) => neg_av_6_31_port, neg_a(30) => 
                           neg_av_6_30_port, neg_a(29) => neg_av_6_29_port, 
                           neg_a(28) => neg_av_6_28_port, neg_a(27) => 
                           neg_av_6_27_port, neg_a(26) => neg_av_6_26_port, 
                           neg_a(25) => neg_av_6_25_port, neg_a(24) => 
                           neg_av_6_24_port, neg_a(23) => neg_av_6_23_port, 
                           neg_a(22) => neg_av_6_22_port, neg_a(21) => 
                           neg_av_6_21_port, neg_a(20) => neg_av_6_20_port, 
                           neg_a(19) => neg_av_6_19_port, neg_a(18) => 
                           neg_av_6_18_port, neg_a(17) => neg_av_6_17_port, 
                           neg_a(16) => neg_av_6_16_port, neg_a(15) => 
                           neg_av_6_15_port, neg_a(14) => neg_av_6_14_port, 
                           neg_a(13) => neg_av_6_13_port, neg_a(12) => 
                           neg_av_6_12_port, neg_a(11) => n_1313, neg_a(10) => 
                           n_1314, neg_a(9) => n_1315, neg_a(8) => n_1316, 
                           neg_a(7) => n_1317, neg_a(6) => n_1318, neg_a(5) => 
                           n_1319, neg_a(4) => n_1320, neg_a(3) => n_1321, 
                           neg_a(2) => n_1322, neg_a(1) => n_1323, neg_a(0) => 
                           n_1324, pos_2a(31) => pos_2av_6_31_port, pos_2a(30) 
                           => pos_2av_6_30_port, pos_2a(29) => 
                           pos_2av_6_29_port, pos_2a(28) => pos_2av_6_28_port, 
                           pos_2a(27) => pos_2av_6_27_port, pos_2a(26) => 
                           pos_2av_6_26_port, pos_2a(25) => pos_2av_6_25_port, 
                           pos_2a(24) => pos_2av_6_24_port, pos_2a(23) => 
                           pos_2av_6_23_port, pos_2a(22) => pos_2av_6_22_port, 
                           pos_2a(21) => pos_2av_6_21_port, pos_2a(20) => 
                           pos_2av_6_20_port, pos_2a(19) => pos_2av_6_19_port, 
                           pos_2a(18) => pos_2av_6_18_port, pos_2a(17) => 
                           pos_2av_6_17_port, pos_2a(16) => pos_2av_6_16_port, 
                           pos_2a(15) => pos_2av_6_15_port, pos_2a(14) => 
                           pos_2av_6_14_port, pos_2a(13) => pos_2av_6_13_port, 
                           pos_2a(12) => n_1325, pos_2a(11) => n_1326, 
                           pos_2a(10) => n_1327, pos_2a(9) => n_1328, pos_2a(8)
                           => n_1329, pos_2a(7) => n_1330, pos_2a(6) => n_1331,
                           pos_2a(5) => n_1332, pos_2a(4) => n_1333, pos_2a(3) 
                           => n_1334, pos_2a(2) => n_1335, pos_2a(1) => n_1336,
                           pos_2a(0) => n_1337, neg_2a(31) => neg_2av_6_31_port
                           , neg_2a(30) => neg_2av_6_30_port, neg_2a(29) => 
                           neg_2av_6_29_port, neg_2a(28) => neg_2av_6_28_port, 
                           neg_2a(27) => neg_2av_6_27_port, neg_2a(26) => 
                           neg_2av_6_26_port, neg_2a(25) => neg_2av_6_25_port, 
                           neg_2a(24) => neg_2av_6_24_port, neg_2a(23) => 
                           neg_2av_6_23_port, neg_2a(22) => neg_2av_6_22_port, 
                           neg_2a(21) => neg_2av_6_21_port, neg_2a(20) => 
                           neg_2av_6_20_port, neg_2a(19) => neg_2av_6_19_port, 
                           neg_2a(18) => neg_2av_6_18_port, neg_2a(17) => 
                           neg_2av_6_17_port, neg_2a(16) => neg_2av_6_16_port, 
                           neg_2a(15) => neg_2av_6_15_port, neg_2a(14) => 
                           neg_2av_6_14_port, neg_2a(13) => neg_2av_6_13_port, 
                           neg_2a(12) => n_1338, neg_2a(11) => n_1339, 
                           neg_2a(10) => n_1340, neg_2a(9) => n_1341, neg_2a(8)
                           => n_1342, neg_2a(7) => n_1343, neg_2a(6) => n_1344,
                           neg_2a(5) => n_1345, neg_2a(4) => n_1346, neg_2a(3) 
                           => n_1347, neg_2a(2) => n_1348, neg_2a(1) => n_1349,
                           neg_2a(0) => n_1350);
   vpn_6 : vp_NBIT32_2 port map( pos_a(31) => pos_av_6_31_port, pos_a(30) => 
                           pos_av_6_30_port, pos_a(29) => pos_av_6_29_port, 
                           pos_a(28) => pos_av_6_28_port, pos_a(27) => 
                           pos_av_6_27_port, pos_a(26) => pos_av_6_26_port, 
                           pos_a(25) => pos_av_6_25_port, pos_a(24) => 
                           pos_av_6_24_port, pos_a(23) => pos_av_6_23_port, 
                           pos_a(22) => pos_av_6_22_port, pos_a(21) => 
                           pos_av_6_21_port, pos_a(20) => pos_av_6_20_port, 
                           pos_a(19) => pos_av_6_19_port, pos_a(18) => 
                           pos_av_6_18_port, pos_a(17) => pos_av_6_17_port, 
                           pos_a(16) => pos_av_6_16_port, pos_a(15) => 
                           pos_av_6_15_port, pos_a(14) => pos_av_6_14_port, 
                           pos_a(13) => pos_av_6_13_port, pos_a(12) => 
                           pos_av_6_12_port, pos_a(11) => pos_av_6_11_port, 
                           pos_a(10) => pos_av_6_10_port, pos_a(9) => 
                           pos_av_6_9_port, pos_a(8) => pos_av_6_8_port, 
                           pos_a(7) => pos_av_6_7_port, pos_a(6) => 
                           pos_av_6_6_port, pos_a(5) => pos_av_6_5_port, 
                           pos_a(4) => pos_av_6_4_port, pos_a(3) => 
                           pos_av_6_3_port, pos_a(2) => pos_av_6_2_port, 
                           pos_a(1) => pos_av_6_1_port, pos_a(0) => 
                           pos_av_6_0_port, neg_a(31) => neg_av_6_31_port, 
                           neg_a(30) => neg_av_6_30_port, neg_a(29) => 
                           neg_av_6_29_port, neg_a(28) => neg_av_6_28_port, 
                           neg_a(27) => neg_av_6_27_port, neg_a(26) => 
                           neg_av_6_26_port, neg_a(25) => neg_av_6_25_port, 
                           neg_a(24) => neg_av_6_24_port, neg_a(23) => 
                           neg_av_6_23_port, neg_a(22) => neg_av_6_22_port, 
                           neg_a(21) => neg_av_6_21_port, neg_a(20) => 
                           neg_av_6_20_port, neg_a(19) => neg_av_6_19_port, 
                           neg_a(18) => neg_av_6_18_port, neg_a(17) => 
                           neg_av_6_17_port, neg_a(16) => neg_av_6_16_port, 
                           neg_a(15) => neg_av_6_15_port, neg_a(14) => 
                           neg_av_6_14_port, neg_a(13) => neg_av_6_13_port, 
                           neg_a(12) => neg_av_6_12_port, neg_a(11) => 
                           neg_av_6_11_port, neg_a(10) => neg_av_6_10_port, 
                           neg_a(9) => neg_av_6_9_port, neg_a(8) => 
                           neg_av_6_8_port, neg_a(7) => neg_av_6_7_port, 
                           neg_a(6) => neg_av_6_6_port, neg_a(5) => 
                           neg_av_6_5_port, neg_a(4) => neg_av_6_4_port, 
                           neg_a(3) => neg_av_6_3_port, neg_a(2) => 
                           neg_av_6_2_port, neg_a(1) => neg_av_6_1_port, 
                           neg_a(0) => neg_av_6_0_port, pos_2a(31) => 
                           pos_2av_6_31_port, pos_2a(30) => pos_2av_6_30_port, 
                           pos_2a(29) => pos_2av_6_29_port, pos_2a(28) => 
                           pos_2av_6_28_port, pos_2a(27) => pos_2av_6_27_port, 
                           pos_2a(26) => pos_2av_6_26_port, pos_2a(25) => 
                           pos_2av_6_25_port, pos_2a(24) => pos_2av_6_24_port, 
                           pos_2a(23) => pos_2av_6_23_port, pos_2a(22) => 
                           pos_2av_6_22_port, pos_2a(21) => pos_2av_6_21_port, 
                           pos_2a(20) => pos_2av_6_20_port, pos_2a(19) => 
                           pos_2av_6_19_port, pos_2a(18) => pos_2av_6_18_port, 
                           pos_2a(17) => pos_2av_6_17_port, pos_2a(16) => 
                           pos_2av_6_16_port, pos_2a(15) => pos_2av_6_15_port, 
                           pos_2a(14) => pos_2av_6_14_port, pos_2a(13) => 
                           pos_2av_6_13_port, pos_2a(12) => pos_2av_6_12_port, 
                           pos_2a(11) => pos_2av_6_11_port, pos_2a(10) => 
                           pos_2av_6_10_port, pos_2a(9) => pos_2av_6_9_port, 
                           pos_2a(8) => pos_2av_6_8_port, pos_2a(7) => 
                           pos_2av_6_7_port, pos_2a(6) => pos_2av_6_6_port, 
                           pos_2a(5) => pos_2av_6_5_port, pos_2a(4) => 
                           pos_2av_6_4_port, pos_2a(3) => pos_2av_6_3_port, 
                           pos_2a(2) => pos_2av_6_2_port, pos_2a(1) => 
                           pos_2av_6_1_port, pos_2a(0) => pos_2av_6_0_port, 
                           neg_2a(31) => neg_2av_6_31_port, neg_2a(30) => 
                           neg_2av_6_30_port, neg_2a(29) => neg_2av_6_29_port, 
                           neg_2a(28) => neg_2av_6_28_port, neg_2a(27) => 
                           neg_2av_6_27_port, neg_2a(26) => neg_2av_6_26_port, 
                           neg_2a(25) => neg_2av_6_25_port, neg_2a(24) => 
                           neg_2av_6_24_port, neg_2a(23) => neg_2av_6_23_port, 
                           neg_2a(22) => neg_2av_6_22_port, neg_2a(21) => 
                           neg_2av_6_21_port, neg_2a(20) => neg_2av_6_20_port, 
                           neg_2a(19) => neg_2av_6_19_port, neg_2a(18) => 
                           neg_2av_6_18_port, neg_2a(17) => neg_2av_6_17_port, 
                           neg_2a(16) => neg_2av_6_16_port, neg_2a(15) => 
                           neg_2av_6_15_port, neg_2a(14) => neg_2av_6_14_port, 
                           neg_2a(13) => neg_2av_6_13_port, neg_2a(12) => 
                           neg_2av_6_12_port, neg_2a(11) => neg_2av_6_11_port, 
                           neg_2a(10) => neg_2av_6_10_port, neg_2a(9) => 
                           neg_2av_6_9_port, neg_2a(8) => neg_2av_6_8_port, 
                           neg_2a(7) => neg_2av_6_7_port, neg_2a(6) => 
                           neg_2av_6_6_port, neg_2a(5) => neg_2av_6_5_port, 
                           neg_2a(4) => neg_2av_6_4_port, neg_2a(3) => 
                           neg_2av_6_3_port, neg_2a(2) => neg_2av_6_2_port, 
                           neg_2a(1) => neg_2av_6_1_port, neg_2a(0) => 
                           neg_2av_6_0_port, sel(2) => b(13), sel(1) => b(12), 
                           sel(0) => b(11), s_out(31) => sum_vector_11_31_port,
                           s_out(30) => sum_vector_11_30_port, s_out(29) => 
                           sum_vector_11_29_port, s_out(28) => 
                           sum_vector_11_28_port, s_out(27) => 
                           sum_vector_11_27_port, s_out(26) => 
                           sum_vector_11_26_port, s_out(25) => 
                           sum_vector_11_25_port, s_out(24) => 
                           sum_vector_11_24_port, s_out(23) => 
                           sum_vector_11_23_port, s_out(22) => 
                           sum_vector_11_22_port, s_out(21) => 
                           sum_vector_11_21_port, s_out(20) => 
                           sum_vector_11_20_port, s_out(19) => 
                           sum_vector_11_19_port, s_out(18) => 
                           sum_vector_11_18_port, s_out(17) => 
                           sum_vector_11_17_port, s_out(16) => 
                           sum_vector_11_16_port, s_out(15) => 
                           sum_vector_11_15_port, s_out(14) => 
                           sum_vector_11_14_port, s_out(13) => 
                           sum_vector_11_13_port, s_out(12) => 
                           sum_vector_11_12_port, s_out(11) => 
                           sum_vector_11_11_port, s_out(10) => 
                           sum_vector_11_10_port, s_out(9) => 
                           sum_vector_11_9_port, s_out(8) => 
                           sum_vector_11_8_port, s_out(7) => 
                           sum_vector_11_7_port, s_out(6) => 
                           sum_vector_11_6_port, s_out(5) => 
                           sum_vector_11_5_port, s_out(4) => 
                           sum_vector_11_4_port, s_out(3) => 
                           sum_vector_11_3_port, s_out(2) => 
                           sum_vector_11_2_port, s_out(1) => 
                           sum_vector_11_1_port, s_out(0) => 
                           sum_vector_11_0_port);
   sumn_6 : rca_signed_NBIT32_2 port map( a(31) => sum_vector_10_31_port, a(30)
                           => sum_vector_10_30_port, a(29) => 
                           sum_vector_10_29_port, a(28) => 
                           sum_vector_10_28_port, a(27) => 
                           sum_vector_10_27_port, a(26) => 
                           sum_vector_10_26_port, a(25) => 
                           sum_vector_10_25_port, a(24) => 
                           sum_vector_10_24_port, a(23) => 
                           sum_vector_10_23_port, a(22) => 
                           sum_vector_10_22_port, a(21) => 
                           sum_vector_10_21_port, a(20) => 
                           sum_vector_10_20_port, a(19) => 
                           sum_vector_10_19_port, a(18) => 
                           sum_vector_10_18_port, a(17) => 
                           sum_vector_10_17_port, a(16) => 
                           sum_vector_10_16_port, a(15) => 
                           sum_vector_10_15_port, a(14) => 
                           sum_vector_10_14_port, a(13) => 
                           sum_vector_10_13_port, a(12) => 
                           sum_vector_10_12_port, a(11) => 
                           sum_vector_10_11_port, a(10) => 
                           sum_vector_10_10_port, a(9) => sum_vector_10_9_port,
                           a(8) => sum_vector_10_8_port, a(7) => 
                           sum_vector_10_7_port, a(6) => sum_vector_10_6_port, 
                           a(5) => sum_vector_10_5_port, a(4) => 
                           sum_vector_10_4_port, a(3) => sum_vector_10_3_port, 
                           a(2) => sum_vector_10_2_port, a(1) => 
                           sum_vector_10_1_port, a(0) => sum_vector_10_0_port, 
                           b(31) => sum_vector_11_31_port, b(30) => 
                           sum_vector_11_30_port, b(29) => 
                           sum_vector_11_29_port, b(28) => 
                           sum_vector_11_28_port, b(27) => 
                           sum_vector_11_27_port, b(26) => 
                           sum_vector_11_26_port, b(25) => 
                           sum_vector_11_25_port, b(24) => 
                           sum_vector_11_24_port, b(23) => 
                           sum_vector_11_23_port, b(22) => 
                           sum_vector_11_22_port, b(21) => 
                           sum_vector_11_21_port, b(20) => 
                           sum_vector_11_20_port, b(19) => 
                           sum_vector_11_19_port, b(18) => 
                           sum_vector_11_18_port, b(17) => 
                           sum_vector_11_17_port, b(16) => 
                           sum_vector_11_16_port, b(15) => 
                           sum_vector_11_15_port, b(14) => 
                           sum_vector_11_14_port, b(13) => 
                           sum_vector_11_13_port, b(12) => 
                           sum_vector_11_12_port, b(11) => 
                           sum_vector_11_11_port, b(10) => 
                           sum_vector_11_10_port, b(9) => sum_vector_11_9_port,
                           b(8) => sum_vector_11_8_port, b(7) => 
                           sum_vector_11_7_port, b(6) => sum_vector_11_6_port, 
                           b(5) => sum_vector_11_5_port, b(4) => 
                           sum_vector_11_4_port, b(3) => sum_vector_11_3_port, 
                           b(2) => sum_vector_11_2_port, b(1) => 
                           sum_vector_11_1_port, b(0) => sum_vector_11_0_port, 
                           c => n_1351, s(31) => sum_vector_12_31_port, s(30) 
                           => sum_vector_12_30_port, s(29) => 
                           sum_vector_12_29_port, s(28) => 
                           sum_vector_12_28_port, s(27) => 
                           sum_vector_12_27_port, s(26) => 
                           sum_vector_12_26_port, s(25) => 
                           sum_vector_12_25_port, s(24) => 
                           sum_vector_12_24_port, s(23) => 
                           sum_vector_12_23_port, s(22) => 
                           sum_vector_12_22_port, s(21) => 
                           sum_vector_12_21_port, s(20) => 
                           sum_vector_12_20_port, s(19) => 
                           sum_vector_12_19_port, s(18) => 
                           sum_vector_12_18_port, s(17) => 
                           sum_vector_12_17_port, s(16) => 
                           sum_vector_12_16_port, s(15) => 
                           sum_vector_12_15_port, s(14) => 
                           sum_vector_12_14_port, s(13) => 
                           sum_vector_12_13_port, s(12) => 
                           sum_vector_12_12_port, s(11) => 
                           sum_vector_12_11_port, s(10) => 
                           sum_vector_12_10_port, s(9) => sum_vector_12_9_port,
                           s(8) => sum_vector_12_8_port, s(7) => 
                           sum_vector_12_7_port, s(6) => sum_vector_12_6_port, 
                           s(5) => sum_vector_12_5_port, s(4) => 
                           sum_vector_12_4_port, s(3) => sum_vector_12_3_port, 
                           s(2) => sum_vector_12_2_port, s(1) => 
                           sum_vector_12_1_port, s(0) => sum_vector_12_0_port);
   shn_7 : shift_NBIT32_SHIFT7 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           pos_a(31) => pos_av_7_31_port, pos_a(30) => 
                           pos_av_7_30_port, pos_a(29) => pos_av_7_29_port, 
                           pos_a(28) => pos_av_7_28_port, pos_a(27) => 
                           pos_av_7_27_port, pos_a(26) => pos_av_7_26_port, 
                           pos_a(25) => pos_av_7_25_port, pos_a(24) => 
                           pos_av_7_24_port, pos_a(23) => pos_av_7_23_port, 
                           pos_a(22) => pos_av_7_22_port, pos_a(21) => 
                           pos_av_7_21_port, pos_a(20) => pos_av_7_20_port, 
                           pos_a(19) => pos_av_7_19_port, pos_a(18) => 
                           pos_av_7_18_port, pos_a(17) => pos_av_7_17_port, 
                           pos_a(16) => pos_av_7_16_port, pos_a(15) => 
                           pos_av_7_15_port, pos_a(14) => pos_av_7_14_port, 
                           pos_a(13) => n_1352, pos_a(12) => n_1353, pos_a(11) 
                           => n_1354, pos_a(10) => n_1355, pos_a(9) => n_1356, 
                           pos_a(8) => n_1357, pos_a(7) => n_1358, pos_a(6) => 
                           n_1359, pos_a(5) => n_1360, pos_a(4) => n_1361, 
                           pos_a(3) => n_1362, pos_a(2) => n_1363, pos_a(1) => 
                           n_1364, pos_a(0) => n_1365, neg_a(31) => 
                           neg_av_7_31_port, neg_a(30) => neg_av_7_30_port, 
                           neg_a(29) => neg_av_7_29_port, neg_a(28) => 
                           neg_av_7_28_port, neg_a(27) => neg_av_7_27_port, 
                           neg_a(26) => neg_av_7_26_port, neg_a(25) => 
                           neg_av_7_25_port, neg_a(24) => neg_av_7_24_port, 
                           neg_a(23) => neg_av_7_23_port, neg_a(22) => 
                           neg_av_7_22_port, neg_a(21) => neg_av_7_21_port, 
                           neg_a(20) => neg_av_7_20_port, neg_a(19) => 
                           neg_av_7_19_port, neg_a(18) => neg_av_7_18_port, 
                           neg_a(17) => neg_av_7_17_port, neg_a(16) => 
                           neg_av_7_16_port, neg_a(15) => neg_av_7_15_port, 
                           neg_a(14) => neg_av_7_14_port, neg_a(13) => n_1366, 
                           neg_a(12) => n_1367, neg_a(11) => n_1368, neg_a(10) 
                           => n_1369, neg_a(9) => n_1370, neg_a(8) => n_1371, 
                           neg_a(7) => n_1372, neg_a(6) => n_1373, neg_a(5) => 
                           n_1374, neg_a(4) => n_1375, neg_a(3) => n_1376, 
                           neg_a(2) => n_1377, neg_a(1) => n_1378, neg_a(0) => 
                           n_1379, pos_2a(31) => pos_2av_7_31_port, pos_2a(30) 
                           => pos_2av_7_30_port, pos_2a(29) => 
                           pos_2av_7_29_port, pos_2a(28) => pos_2av_7_28_port, 
                           pos_2a(27) => pos_2av_7_27_port, pos_2a(26) => 
                           pos_2av_7_26_port, pos_2a(25) => pos_2av_7_25_port, 
                           pos_2a(24) => pos_2av_7_24_port, pos_2a(23) => 
                           pos_2av_7_23_port, pos_2a(22) => pos_2av_7_22_port, 
                           pos_2a(21) => pos_2av_7_21_port, pos_2a(20) => 
                           pos_2av_7_20_port, pos_2a(19) => pos_2av_7_19_port, 
                           pos_2a(18) => pos_2av_7_18_port, pos_2a(17) => 
                           pos_2av_7_17_port, pos_2a(16) => pos_2av_7_16_port, 
                           pos_2a(15) => pos_2av_7_15_port, pos_2a(14) => 
                           n_1380, pos_2a(13) => n_1381, pos_2a(12) => n_1382, 
                           pos_2a(11) => n_1383, pos_2a(10) => n_1384, 
                           pos_2a(9) => n_1385, pos_2a(8) => n_1386, pos_2a(7) 
                           => n_1387, pos_2a(6) => n_1388, pos_2a(5) => n_1389,
                           pos_2a(4) => n_1390, pos_2a(3) => n_1391, pos_2a(2) 
                           => n_1392, pos_2a(1) => n_1393, pos_2a(0) => n_1394,
                           neg_2a(31) => neg_2av_7_31_port, neg_2a(30) => 
                           neg_2av_7_30_port, neg_2a(29) => neg_2av_7_29_port, 
                           neg_2a(28) => neg_2av_7_28_port, neg_2a(27) => 
                           neg_2av_7_27_port, neg_2a(26) => neg_2av_7_26_port, 
                           neg_2a(25) => neg_2av_7_25_port, neg_2a(24) => 
                           neg_2av_7_24_port, neg_2a(23) => neg_2av_7_23_port, 
                           neg_2a(22) => neg_2av_7_22_port, neg_2a(21) => 
                           neg_2av_7_21_port, neg_2a(20) => neg_2av_7_20_port, 
                           neg_2a(19) => neg_2av_7_19_port, neg_2a(18) => 
                           neg_2av_7_18_port, neg_2a(17) => neg_2av_7_17_port, 
                           neg_2a(16) => neg_2av_7_16_port, neg_2a(15) => 
                           neg_2av_7_15_port, neg_2a(14) => n_1395, neg_2a(13) 
                           => n_1396, neg_2a(12) => n_1397, neg_2a(11) => 
                           n_1398, neg_2a(10) => n_1399, neg_2a(9) => n_1400, 
                           neg_2a(8) => n_1401, neg_2a(7) => n_1402, neg_2a(6) 
                           => n_1403, neg_2a(5) => n_1404, neg_2a(4) => n_1405,
                           neg_2a(3) => n_1406, neg_2a(2) => n_1407, neg_2a(1) 
                           => n_1408, neg_2a(0) => n_1409);
   vpn_7 : vp_NBIT32_1 port map( pos_a(31) => pos_av_7_31_port, pos_a(30) => 
                           pos_av_7_30_port, pos_a(29) => pos_av_7_29_port, 
                           pos_a(28) => pos_av_7_28_port, pos_a(27) => 
                           pos_av_7_27_port, pos_a(26) => pos_av_7_26_port, 
                           pos_a(25) => pos_av_7_25_port, pos_a(24) => 
                           pos_av_7_24_port, pos_a(23) => pos_av_7_23_port, 
                           pos_a(22) => pos_av_7_22_port, pos_a(21) => 
                           pos_av_7_21_port, pos_a(20) => pos_av_7_20_port, 
                           pos_a(19) => pos_av_7_19_port, pos_a(18) => 
                           pos_av_7_18_port, pos_a(17) => pos_av_7_17_port, 
                           pos_a(16) => pos_av_7_16_port, pos_a(15) => 
                           pos_av_7_15_port, pos_a(14) => pos_av_7_14_port, 
                           pos_a(13) => pos_av_7_13_port, pos_a(12) => 
                           pos_av_7_12_port, pos_a(11) => pos_av_7_11_port, 
                           pos_a(10) => pos_av_7_10_port, pos_a(9) => 
                           pos_av_7_9_port, pos_a(8) => pos_av_7_8_port, 
                           pos_a(7) => pos_av_7_7_port, pos_a(6) => 
                           pos_av_7_6_port, pos_a(5) => pos_av_7_5_port, 
                           pos_a(4) => pos_av_7_4_port, pos_a(3) => 
                           pos_av_7_3_port, pos_a(2) => pos_av_7_2_port, 
                           pos_a(1) => pos_av_7_1_port, pos_a(0) => 
                           pos_av_7_0_port, neg_a(31) => neg_av_7_31_port, 
                           neg_a(30) => neg_av_7_30_port, neg_a(29) => 
                           neg_av_7_29_port, neg_a(28) => neg_av_7_28_port, 
                           neg_a(27) => neg_av_7_27_port, neg_a(26) => 
                           neg_av_7_26_port, neg_a(25) => neg_av_7_25_port, 
                           neg_a(24) => neg_av_7_24_port, neg_a(23) => 
                           neg_av_7_23_port, neg_a(22) => neg_av_7_22_port, 
                           neg_a(21) => neg_av_7_21_port, neg_a(20) => 
                           neg_av_7_20_port, neg_a(19) => neg_av_7_19_port, 
                           neg_a(18) => neg_av_7_18_port, neg_a(17) => 
                           neg_av_7_17_port, neg_a(16) => neg_av_7_16_port, 
                           neg_a(15) => neg_av_7_15_port, neg_a(14) => 
                           neg_av_7_14_port, neg_a(13) => neg_av_7_13_port, 
                           neg_a(12) => neg_av_7_12_port, neg_a(11) => 
                           neg_av_7_11_port, neg_a(10) => neg_av_7_10_port, 
                           neg_a(9) => neg_av_7_9_port, neg_a(8) => 
                           neg_av_7_8_port, neg_a(7) => neg_av_7_7_port, 
                           neg_a(6) => neg_av_7_6_port, neg_a(5) => 
                           neg_av_7_5_port, neg_a(4) => neg_av_7_4_port, 
                           neg_a(3) => neg_av_7_3_port, neg_a(2) => 
                           neg_av_7_2_port, neg_a(1) => neg_av_7_1_port, 
                           neg_a(0) => neg_av_7_0_port, pos_2a(31) => 
                           pos_2av_7_31_port, pos_2a(30) => pos_2av_7_30_port, 
                           pos_2a(29) => pos_2av_7_29_port, pos_2a(28) => 
                           pos_2av_7_28_port, pos_2a(27) => pos_2av_7_27_port, 
                           pos_2a(26) => pos_2av_7_26_port, pos_2a(25) => 
                           pos_2av_7_25_port, pos_2a(24) => pos_2av_7_24_port, 
                           pos_2a(23) => pos_2av_7_23_port, pos_2a(22) => 
                           pos_2av_7_22_port, pos_2a(21) => pos_2av_7_21_port, 
                           pos_2a(20) => pos_2av_7_20_port, pos_2a(19) => 
                           pos_2av_7_19_port, pos_2a(18) => pos_2av_7_18_port, 
                           pos_2a(17) => pos_2av_7_17_port, pos_2a(16) => 
                           pos_2av_7_16_port, pos_2a(15) => pos_2av_7_15_port, 
                           pos_2a(14) => pos_2av_7_14_port, pos_2a(13) => 
                           pos_2av_7_13_port, pos_2a(12) => pos_2av_7_12_port, 
                           pos_2a(11) => pos_2av_7_11_port, pos_2a(10) => 
                           pos_2av_7_10_port, pos_2a(9) => pos_2av_7_9_port, 
                           pos_2a(8) => pos_2av_7_8_port, pos_2a(7) => 
                           pos_2av_7_7_port, pos_2a(6) => pos_2av_7_6_port, 
                           pos_2a(5) => pos_2av_7_5_port, pos_2a(4) => 
                           pos_2av_7_4_port, pos_2a(3) => pos_2av_7_3_port, 
                           pos_2a(2) => pos_2av_7_2_port, pos_2a(1) => 
                           pos_2av_7_1_port, pos_2a(0) => pos_2av_7_0_port, 
                           neg_2a(31) => neg_2av_7_31_port, neg_2a(30) => 
                           neg_2av_7_30_port, neg_2a(29) => neg_2av_7_29_port, 
                           neg_2a(28) => neg_2av_7_28_port, neg_2a(27) => 
                           neg_2av_7_27_port, neg_2a(26) => neg_2av_7_26_port, 
                           neg_2a(25) => neg_2av_7_25_port, neg_2a(24) => 
                           neg_2av_7_24_port, neg_2a(23) => neg_2av_7_23_port, 
                           neg_2a(22) => neg_2av_7_22_port, neg_2a(21) => 
                           neg_2av_7_21_port, neg_2a(20) => neg_2av_7_20_port, 
                           neg_2a(19) => neg_2av_7_19_port, neg_2a(18) => 
                           neg_2av_7_18_port, neg_2a(17) => neg_2av_7_17_port, 
                           neg_2a(16) => neg_2av_7_16_port, neg_2a(15) => 
                           neg_2av_7_15_port, neg_2a(14) => neg_2av_7_14_port, 
                           neg_2a(13) => neg_2av_7_13_port, neg_2a(12) => 
                           neg_2av_7_12_port, neg_2a(11) => neg_2av_7_11_port, 
                           neg_2a(10) => neg_2av_7_10_port, neg_2a(9) => 
                           neg_2av_7_9_port, neg_2a(8) => neg_2av_7_8_port, 
                           neg_2a(7) => neg_2av_7_7_port, neg_2a(6) => 
                           neg_2av_7_6_port, neg_2a(5) => neg_2av_7_5_port, 
                           neg_2a(4) => neg_2av_7_4_port, neg_2a(3) => 
                           neg_2av_7_3_port, neg_2a(2) => neg_2av_7_2_port, 
                           neg_2a(1) => neg_2av_7_1_port, neg_2a(0) => 
                           neg_2av_7_0_port, sel(2) => b(15), sel(1) => b(14), 
                           sel(0) => b(13), s_out(31) => sum_vector_13_31_port,
                           s_out(30) => sum_vector_13_30_port, s_out(29) => 
                           sum_vector_13_29_port, s_out(28) => 
                           sum_vector_13_28_port, s_out(27) => 
                           sum_vector_13_27_port, s_out(26) => 
                           sum_vector_13_26_port, s_out(25) => 
                           sum_vector_13_25_port, s_out(24) => 
                           sum_vector_13_24_port, s_out(23) => 
                           sum_vector_13_23_port, s_out(22) => 
                           sum_vector_13_22_port, s_out(21) => 
                           sum_vector_13_21_port, s_out(20) => 
                           sum_vector_13_20_port, s_out(19) => 
                           sum_vector_13_19_port, s_out(18) => 
                           sum_vector_13_18_port, s_out(17) => 
                           sum_vector_13_17_port, s_out(16) => 
                           sum_vector_13_16_port, s_out(15) => 
                           sum_vector_13_15_port, s_out(14) => 
                           sum_vector_13_14_port, s_out(13) => 
                           sum_vector_13_13_port, s_out(12) => 
                           sum_vector_13_12_port, s_out(11) => 
                           sum_vector_13_11_port, s_out(10) => 
                           sum_vector_13_10_port, s_out(9) => 
                           sum_vector_13_9_port, s_out(8) => 
                           sum_vector_13_8_port, s_out(7) => 
                           sum_vector_13_7_port, s_out(6) => 
                           sum_vector_13_6_port, s_out(5) => 
                           sum_vector_13_5_port, s_out(4) => 
                           sum_vector_13_4_port, s_out(3) => 
                           sum_vector_13_3_port, s_out(2) => 
                           sum_vector_13_2_port, s_out(1) => 
                           sum_vector_13_1_port, s_out(0) => 
                           sum_vector_13_0_port);
   sumn_7 : rca_signed_NBIT32_1 port map( a(31) => sum_vector_12_31_port, a(30)
                           => sum_vector_12_30_port, a(29) => 
                           sum_vector_12_29_port, a(28) => 
                           sum_vector_12_28_port, a(27) => 
                           sum_vector_12_27_port, a(26) => 
                           sum_vector_12_26_port, a(25) => 
                           sum_vector_12_25_port, a(24) => 
                           sum_vector_12_24_port, a(23) => 
                           sum_vector_12_23_port, a(22) => 
                           sum_vector_12_22_port, a(21) => 
                           sum_vector_12_21_port, a(20) => 
                           sum_vector_12_20_port, a(19) => 
                           sum_vector_12_19_port, a(18) => 
                           sum_vector_12_18_port, a(17) => 
                           sum_vector_12_17_port, a(16) => 
                           sum_vector_12_16_port, a(15) => 
                           sum_vector_12_15_port, a(14) => 
                           sum_vector_12_14_port, a(13) => 
                           sum_vector_12_13_port, a(12) => 
                           sum_vector_12_12_port, a(11) => 
                           sum_vector_12_11_port, a(10) => 
                           sum_vector_12_10_port, a(9) => sum_vector_12_9_port,
                           a(8) => sum_vector_12_8_port, a(7) => 
                           sum_vector_12_7_port, a(6) => sum_vector_12_6_port, 
                           a(5) => sum_vector_12_5_port, a(4) => 
                           sum_vector_12_4_port, a(3) => sum_vector_12_3_port, 
                           a(2) => sum_vector_12_2_port, a(1) => 
                           sum_vector_12_1_port, a(0) => sum_vector_12_0_port, 
                           b(31) => sum_vector_13_31_port, b(30) => 
                           sum_vector_13_30_port, b(29) => 
                           sum_vector_13_29_port, b(28) => 
                           sum_vector_13_28_port, b(27) => 
                           sum_vector_13_27_port, b(26) => 
                           sum_vector_13_26_port, b(25) => 
                           sum_vector_13_25_port, b(24) => 
                           sum_vector_13_24_port, b(23) => 
                           sum_vector_13_23_port, b(22) => 
                           sum_vector_13_22_port, b(21) => 
                           sum_vector_13_21_port, b(20) => 
                           sum_vector_13_20_port, b(19) => 
                           sum_vector_13_19_port, b(18) => 
                           sum_vector_13_18_port, b(17) => 
                           sum_vector_13_17_port, b(16) => 
                           sum_vector_13_16_port, b(15) => 
                           sum_vector_13_15_port, b(14) => 
                           sum_vector_13_14_port, b(13) => 
                           sum_vector_13_13_port, b(12) => 
                           sum_vector_13_12_port, b(11) => 
                           sum_vector_13_11_port, b(10) => 
                           sum_vector_13_10_port, b(9) => sum_vector_13_9_port,
                           b(8) => sum_vector_13_8_port, b(7) => 
                           sum_vector_13_7_port, b(6) => sum_vector_13_6_port, 
                           b(5) => sum_vector_13_5_port, b(4) => 
                           sum_vector_13_4_port, b(3) => sum_vector_13_3_port, 
                           b(2) => sum_vector_13_2_port, b(1) => 
                           sum_vector_13_1_port, b(0) => sum_vector_13_0_port, 
                           c => n_1410, s(31) => mul(31), s(30) => mul(30), 
                           s(29) => mul(29), s(28) => mul(28), s(27) => mul(27)
                           , s(26) => mul(26), s(25) => mul(25), s(24) => 
                           mul(24), s(23) => mul(23), s(22) => mul(22), s(21) 
                           => mul(21), s(20) => mul(20), s(19) => mul(19), 
                           s(18) => mul(18), s(17) => mul(17), s(16) => mul(16)
                           , s(15) => mul(15), s(14) => mul(14), s(13) => 
                           mul(13), s(12) => mul(12), s(11) => mul(11), s(10) 
                           => mul(10), s(9) => mul(9), s(8) => mul(8), s(7) => 
                           mul(7), s(6) => mul(6), s(5) => mul(5), s(4) => 
                           mul(4), s(3) => mul(3), s(2) => mul(2), s(1) => 
                           mul(1), s(0) => mul(0));
   neg_2av_7_0_port <= '0';
   neg_2av_7_1_port <= '0';
   neg_2av_7_2_port <= '0';
   neg_2av_7_3_port <= '0';
   neg_2av_7_4_port <= '0';
   neg_2av_7_5_port <= '0';
   neg_2av_7_6_port <= '0';
   neg_2av_7_7_port <= '0';
   neg_2av_7_8_port <= '0';
   neg_2av_7_9_port <= '0';
   neg_2av_7_10_port <= '0';
   neg_2av_7_11_port <= '0';
   neg_2av_7_12_port <= '0';
   neg_2av_7_13_port <= '0';
   neg_2av_7_14_port <= '0';
   pos_2av_7_0_port <= '0';
   pos_2av_7_1_port <= '0';
   pos_2av_7_2_port <= '0';
   pos_2av_7_3_port <= '0';
   pos_2av_7_4_port <= '0';
   pos_2av_7_5_port <= '0';
   pos_2av_7_6_port <= '0';
   pos_2av_7_7_port <= '0';
   pos_2av_7_8_port <= '0';
   pos_2av_7_9_port <= '0';
   pos_2av_7_10_port <= '0';
   pos_2av_7_11_port <= '0';
   pos_2av_7_12_port <= '0';
   pos_2av_7_13_port <= '0';
   pos_2av_7_14_port <= '0';
   neg_av_7_0_port <= '0';
   neg_av_7_1_port <= '0';
   neg_av_7_2_port <= '0';
   neg_av_7_3_port <= '0';
   neg_av_7_4_port <= '0';
   neg_av_7_5_port <= '0';
   neg_av_7_6_port <= '0';
   neg_av_7_7_port <= '0';
   neg_av_7_8_port <= '0';
   neg_av_7_9_port <= '0';
   neg_av_7_10_port <= '0';
   neg_av_7_11_port <= '0';
   neg_av_7_12_port <= '0';
   neg_av_7_13_port <= '0';
   pos_av_7_0_port <= '0';
   pos_av_7_1_port <= '0';
   pos_av_7_2_port <= '0';
   pos_av_7_3_port <= '0';
   pos_av_7_4_port <= '0';
   pos_av_7_5_port <= '0';
   pos_av_7_6_port <= '0';
   pos_av_7_7_port <= '0';
   pos_av_7_8_port <= '0';
   pos_av_7_9_port <= '0';
   pos_av_7_10_port <= '0';
   pos_av_7_11_port <= '0';
   pos_av_7_12_port <= '0';
   pos_av_7_13_port <= '0';
   neg_2av_6_0_port <= '0';
   neg_2av_6_1_port <= '0';
   neg_2av_6_2_port <= '0';
   neg_2av_6_3_port <= '0';
   neg_2av_6_4_port <= '0';
   neg_2av_6_5_port <= '0';
   neg_2av_6_6_port <= '0';
   neg_2av_6_7_port <= '0';
   neg_2av_6_8_port <= '0';
   neg_2av_6_9_port <= '0';
   neg_2av_6_10_port <= '0';
   neg_2av_6_11_port <= '0';
   neg_2av_6_12_port <= '0';
   pos_2av_6_0_port <= '0';
   pos_2av_6_1_port <= '0';
   pos_2av_6_2_port <= '0';
   pos_2av_6_3_port <= '0';
   pos_2av_6_4_port <= '0';
   pos_2av_6_5_port <= '0';
   pos_2av_6_6_port <= '0';
   pos_2av_6_7_port <= '0';
   pos_2av_6_8_port <= '0';
   pos_2av_6_9_port <= '0';
   pos_2av_6_10_port <= '0';
   pos_2av_6_11_port <= '0';
   pos_2av_6_12_port <= '0';
   neg_av_6_0_port <= '0';
   neg_av_6_1_port <= '0';
   neg_av_6_2_port <= '0';
   neg_av_6_3_port <= '0';
   neg_av_6_4_port <= '0';
   neg_av_6_5_port <= '0';
   neg_av_6_6_port <= '0';
   neg_av_6_7_port <= '0';
   neg_av_6_8_port <= '0';
   neg_av_6_9_port <= '0';
   neg_av_6_10_port <= '0';
   neg_av_6_11_port <= '0';
   pos_av_6_0_port <= '0';
   pos_av_6_1_port <= '0';
   pos_av_6_2_port <= '0';
   pos_av_6_3_port <= '0';
   pos_av_6_4_port <= '0';
   pos_av_6_5_port <= '0';
   pos_av_6_6_port <= '0';
   pos_av_6_7_port <= '0';
   pos_av_6_8_port <= '0';
   pos_av_6_9_port <= '0';
   pos_av_6_10_port <= '0';
   pos_av_6_11_port <= '0';
   neg_2av_5_0_port <= '0';
   neg_2av_5_1_port <= '0';
   neg_2av_5_2_port <= '0';
   neg_2av_5_3_port <= '0';
   neg_2av_5_4_port <= '0';
   neg_2av_5_5_port <= '0';
   neg_2av_5_6_port <= '0';
   neg_2av_5_7_port <= '0';
   neg_2av_5_8_port <= '0';
   neg_2av_5_9_port <= '0';
   neg_2av_5_10_port <= '0';
   pos_2av_5_0_port <= '0';
   pos_2av_5_1_port <= '0';
   pos_2av_5_2_port <= '0';
   pos_2av_5_3_port <= '0';
   pos_2av_5_4_port <= '0';
   pos_2av_5_5_port <= '0';
   pos_2av_5_6_port <= '0';
   pos_2av_5_7_port <= '0';
   pos_2av_5_8_port <= '0';
   pos_2av_5_9_port <= '0';
   pos_2av_5_10_port <= '0';
   neg_av_5_0_port <= '0';
   neg_av_5_1_port <= '0';
   neg_av_5_2_port <= '0';
   neg_av_5_3_port <= '0';
   neg_av_5_4_port <= '0';
   neg_av_5_5_port <= '0';
   neg_av_5_6_port <= '0';
   neg_av_5_7_port <= '0';
   neg_av_5_8_port <= '0';
   neg_av_5_9_port <= '0';
   pos_av_5_0_port <= '0';
   pos_av_5_1_port <= '0';
   pos_av_5_2_port <= '0';
   pos_av_5_3_port <= '0';
   pos_av_5_4_port <= '0';
   pos_av_5_5_port <= '0';
   pos_av_5_6_port <= '0';
   pos_av_5_7_port <= '0';
   pos_av_5_8_port <= '0';
   pos_av_5_9_port <= '0';
   neg_2av_4_0_port <= '0';
   neg_2av_4_1_port <= '0';
   neg_2av_4_2_port <= '0';
   neg_2av_4_3_port <= '0';
   neg_2av_4_4_port <= '0';
   neg_2av_4_5_port <= '0';
   neg_2av_4_6_port <= '0';
   neg_2av_4_7_port <= '0';
   neg_2av_4_8_port <= '0';
   pos_2av_4_0_port <= '0';
   pos_2av_4_1_port <= '0';
   pos_2av_4_2_port <= '0';
   pos_2av_4_3_port <= '0';
   pos_2av_4_4_port <= '0';
   pos_2av_4_5_port <= '0';
   pos_2av_4_6_port <= '0';
   pos_2av_4_7_port <= '0';
   pos_2av_4_8_port <= '0';
   neg_av_4_0_port <= '0';
   neg_av_4_1_port <= '0';
   neg_av_4_2_port <= '0';
   neg_av_4_3_port <= '0';
   neg_av_4_4_port <= '0';
   neg_av_4_5_port <= '0';
   neg_av_4_6_port <= '0';
   neg_av_4_7_port <= '0';
   pos_av_4_0_port <= '0';
   pos_av_4_1_port <= '0';
   pos_av_4_2_port <= '0';
   pos_av_4_3_port <= '0';
   pos_av_4_4_port <= '0';
   pos_av_4_5_port <= '0';
   pos_av_4_6_port <= '0';
   pos_av_4_7_port <= '0';
   neg_2av_3_0_port <= '0';
   neg_2av_3_1_port <= '0';
   neg_2av_3_2_port <= '0';
   neg_2av_3_3_port <= '0';
   neg_2av_3_4_port <= '0';
   neg_2av_3_5_port <= '0';
   neg_2av_3_6_port <= '0';
   pos_2av_3_0_port <= '0';
   pos_2av_3_1_port <= '0';
   pos_2av_3_2_port <= '0';
   pos_2av_3_3_port <= '0';
   pos_2av_3_4_port <= '0';
   pos_2av_3_5_port <= '0';
   pos_2av_3_6_port <= '0';
   neg_av_3_0_port <= '0';
   neg_av_3_1_port <= '0';
   neg_av_3_2_port <= '0';
   neg_av_3_3_port <= '0';
   neg_av_3_4_port <= '0';
   neg_av_3_5_port <= '0';
   pos_av_3_0_port <= '0';
   pos_av_3_1_port <= '0';
   pos_av_3_2_port <= '0';
   pos_av_3_3_port <= '0';
   pos_av_3_4_port <= '0';
   pos_av_3_5_port <= '0';
   neg_2av_2_0_port <= '0';
   neg_2av_2_1_port <= '0';
   neg_2av_2_2_port <= '0';
   neg_2av_2_3_port <= '0';
   neg_2av_2_4_port <= '0';
   pos_2av_2_0_port <= '0';
   pos_2av_2_1_port <= '0';
   pos_2av_2_2_port <= '0';
   pos_2av_2_3_port <= '0';
   pos_2av_2_4_port <= '0';
   neg_av_2_0_port <= '0';
   neg_av_2_1_port <= '0';
   neg_av_2_2_port <= '0';
   neg_av_2_3_port <= '0';
   pos_av_2_0_port <= '0';
   pos_av_2_1_port <= '0';
   pos_av_2_2_port <= '0';
   pos_av_2_3_port <= '0';
   neg_2av_1_0_port <= '0';
   neg_2av_1_1_port <= '0';
   neg_2av_1_2_port <= '0';
   pos_2av_1_0_port <= '0';
   pos_2av_1_1_port <= '0';
   pos_2av_1_2_port <= '0';
   neg_av_1_0_port <= '0';
   neg_av_1_1_port <= '0';
   pos_av_1_0_port <= '0';
   pos_av_1_1_port <= '0';
   neg_2av_0_0_port <= '0';
   pos_2av_0_0_port <= '0';

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity sparse_tree_adder_n_bit32 is

   port( operand_1, operand_2 : in std_logic_vector (31 downto 0);  carry_in : 
         in std_logic;  sum : out std_logic_vector (31 downto 0);  carry_out, 
         overflow : out std_logic);

end sparse_tree_adder_n_bit32;

architecture SYN_specification of sparse_tree_adder_n_bit32 is

   component carry_select_adder_n_bit4_1
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component carry_select_adder_n_bit4_2
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component carry_select_adder_n_bit4_3
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component carry_select_adder_n_bit4_4
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component carry_select_adder_n_bit4_5
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component carry_select_adder_n_bit4_6
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component carry_select_adder_n_bit4_7
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component carry_select_adder_n_bit4_0
      port( operand_1, operand_2 : in std_logic_vector (3 downto 0);  carry_in 
            : in std_logic;  sum : out std_logic_vector (3 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component sparse_tree_carry_generator_n_bit32
      port( operand_1, operand_2 : in std_logic_vector (31 downto 0);  carry_in
            : in std_logic;  carry_out : out std_logic_vector (7 downto 0));
   end component;
   
   signal carries_7_port, carries_6_port, carries_5_port, carries_4_port, 
      carries_3_port, carries_2_port, carries_1_port, n_1411, n_1412, n_1413, 
      n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, 
      n_1423, n_1424, n_1425 : std_logic;

begin
   
   carrygen : sparse_tree_carry_generator_n_bit32 port map( operand_1(31) => 
                           operand_1(31), operand_1(30) => operand_1(30), 
                           operand_1(29) => operand_1(29), operand_1(28) => 
                           operand_1(28), operand_1(27) => operand_1(27), 
                           operand_1(26) => operand_1(26), operand_1(25) => 
                           operand_1(25), operand_1(24) => operand_1(24), 
                           operand_1(23) => operand_1(23), operand_1(22) => 
                           operand_1(22), operand_1(21) => operand_1(21), 
                           operand_1(20) => operand_1(20), operand_1(19) => 
                           operand_1(19), operand_1(18) => operand_1(18), 
                           operand_1(17) => operand_1(17), operand_1(16) => 
                           operand_1(16), operand_1(15) => operand_1(15), 
                           operand_1(14) => operand_1(14), operand_1(13) => 
                           operand_1(13), operand_1(12) => operand_1(12), 
                           operand_1(11) => operand_1(11), operand_1(10) => 
                           operand_1(10), operand_1(9) => operand_1(9), 
                           operand_1(8) => operand_1(8), operand_1(7) => 
                           operand_1(7), operand_1(6) => operand_1(6), 
                           operand_1(5) => operand_1(5), operand_1(4) => 
                           operand_1(4), operand_1(3) => operand_1(3), 
                           operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(31) => operand_2(31), operand_2(30) => 
                           operand_2(30), operand_2(29) => operand_2(29), 
                           operand_2(28) => operand_2(28), operand_2(27) => 
                           operand_2(27), operand_2(26) => operand_2(26), 
                           operand_2(25) => operand_2(25), operand_2(24) => 
                           operand_2(24), operand_2(23) => operand_2(23), 
                           operand_2(22) => operand_2(22), operand_2(21) => 
                           operand_2(21), operand_2(20) => operand_2(20), 
                           operand_2(19) => operand_2(19), operand_2(18) => 
                           operand_2(18), operand_2(17) => operand_2(17), 
                           operand_2(16) => operand_2(16), operand_2(15) => 
                           operand_2(15), operand_2(14) => operand_2(14), 
                           operand_2(13) => operand_2(13), operand_2(12) => 
                           operand_2(12), operand_2(11) => operand_2(11), 
                           operand_2(10) => operand_2(10), operand_2(9) => 
                           operand_2(9), operand_2(8) => operand_2(8), 
                           operand_2(7) => operand_2(7), operand_2(6) => 
                           operand_2(6), operand_2(5) => operand_2(5), 
                           operand_2(4) => operand_2(4), operand_2(3) => 
                           operand_2(3), operand_2(2) => operand_2(2), 
                           operand_2(1) => operand_2(1), operand_2(0) => 
                           operand_2(0), carry_in => carry_in, carry_out(7) => 
                           carry_out, carry_out(6) => carries_7_port, 
                           carry_out(5) => carries_6_port, carry_out(4) => 
                           carries_5_port, carry_out(3) => carries_4_port, 
                           carry_out(2) => carries_3_port, carry_out(1) => 
                           carries_2_port, carry_out(0) => carries_1_port);
   adder_0 : carry_select_adder_n_bit4_0 port map( operand_1(3) => operand_1(3)
                           , operand_1(2) => operand_1(2), operand_1(1) => 
                           operand_1(1), operand_1(0) => operand_1(0), 
                           operand_2(3) => operand_2(3), operand_2(2) => 
                           operand_2(2), operand_2(1) => operand_2(1), 
                           operand_2(0) => operand_2(0), carry_in => carry_in, 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0), carry_out => n_1411, overflow =>
                           n_1412);
   adder_1 : carry_select_adder_n_bit4_7 port map( operand_1(3) => operand_1(7)
                           , operand_1(2) => operand_1(6), operand_1(1) => 
                           operand_1(5), operand_1(0) => operand_1(4), 
                           operand_2(3) => operand_2(7), operand_2(2) => 
                           operand_2(6), operand_2(1) => operand_2(5), 
                           operand_2(0) => operand_2(4), carry_in => 
                           carries_1_port, sum(3) => sum(7), sum(2) => sum(6), 
                           sum(1) => sum(5), sum(0) => sum(4), carry_out => 
                           n_1413, overflow => n_1414);
   adder_2 : carry_select_adder_n_bit4_6 port map( operand_1(3) => 
                           operand_1(11), operand_1(2) => operand_1(10), 
                           operand_1(1) => operand_1(9), operand_1(0) => 
                           operand_1(8), operand_2(3) => operand_2(11), 
                           operand_2(2) => operand_2(10), operand_2(1) => 
                           operand_2(9), operand_2(0) => operand_2(8), carry_in
                           => carries_2_port, sum(3) => sum(11), sum(2) => 
                           sum(10), sum(1) => sum(9), sum(0) => sum(8), 
                           carry_out => n_1415, overflow => n_1416);
   adder_3 : carry_select_adder_n_bit4_5 port map( operand_1(3) => 
                           operand_1(15), operand_1(2) => operand_1(14), 
                           operand_1(1) => operand_1(13), operand_1(0) => 
                           operand_1(12), operand_2(3) => operand_2(15), 
                           operand_2(2) => operand_2(14), operand_2(1) => 
                           operand_2(13), operand_2(0) => operand_2(12), 
                           carry_in => carries_3_port, sum(3) => sum(15), 
                           sum(2) => sum(14), sum(1) => sum(13), sum(0) => 
                           sum(12), carry_out => n_1417, overflow => n_1418);
   adder_4 : carry_select_adder_n_bit4_4 port map( operand_1(3) => 
                           operand_1(19), operand_1(2) => operand_1(18), 
                           operand_1(1) => operand_1(17), operand_1(0) => 
                           operand_1(16), operand_2(3) => operand_2(19), 
                           operand_2(2) => operand_2(18), operand_2(1) => 
                           operand_2(17), operand_2(0) => operand_2(16), 
                           carry_in => carries_4_port, sum(3) => sum(19), 
                           sum(2) => sum(18), sum(1) => sum(17), sum(0) => 
                           sum(16), carry_out => n_1419, overflow => n_1420);
   adder_5 : carry_select_adder_n_bit4_3 port map( operand_1(3) => 
                           operand_1(23), operand_1(2) => operand_1(22), 
                           operand_1(1) => operand_1(21), operand_1(0) => 
                           operand_1(20), operand_2(3) => operand_2(23), 
                           operand_2(2) => operand_2(22), operand_2(1) => 
                           operand_2(21), operand_2(0) => operand_2(20), 
                           carry_in => carries_5_port, sum(3) => sum(23), 
                           sum(2) => sum(22), sum(1) => sum(21), sum(0) => 
                           sum(20), carry_out => n_1421, overflow => n_1422);
   adder_6 : carry_select_adder_n_bit4_2 port map( operand_1(3) => 
                           operand_1(27), operand_1(2) => operand_1(26), 
                           operand_1(1) => operand_1(25), operand_1(0) => 
                           operand_1(24), operand_2(3) => operand_2(27), 
                           operand_2(2) => operand_2(26), operand_2(1) => 
                           operand_2(25), operand_2(0) => operand_2(24), 
                           carry_in => carries_6_port, sum(3) => sum(27), 
                           sum(2) => sum(26), sum(1) => sum(25), sum(0) => 
                           sum(24), carry_out => n_1423, overflow => n_1424);
   adder_7 : carry_select_adder_n_bit4_1 port map( operand_1(3) => 
                           operand_1(31), operand_1(2) => operand_1(30), 
                           operand_1(1) => operand_1(29), operand_1(0) => 
                           operand_1(28), operand_2(3) => operand_2(31), 
                           operand_2(2) => operand_2(30), operand_2(1) => 
                           operand_2(29), operand_2(0) => operand_2(28), 
                           carry_in => carries_7_port, sum(3) => sum(31), 
                           sum(2) => sum(30), sum(1) => sum(29), sum(0) => 
                           sum(28), carry_out => n_1425, overflow => overflow);

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity shifter_wrapper_nbit32 is

   port( r1, r2 : in std_logic_vector (31 downto 0);  conf : in 
         std_logic_vector (1 downto 0);  en_shifter : in std_logic;  
         shifted_out : out std_logic_vector (31 downto 0));

end shifter_wrapper_nbit32;

architecture SYN_behavioral of shifter_wrapper_nbit32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shifter_nbit32
      port( r1, r2 : in std_logic_vector (31 downto 0);  conf : in 
            std_logic_vector (1 downto 0);  shifted_out : out std_logic_vector 
            (31 downto 0));
   end component;
   
   signal shifted_out_i_31_port, shifted_out_i_30_port, shifted_out_i_29_port, 
      shifted_out_i_28_port, shifted_out_i_27_port, shifted_out_i_26_port, 
      shifted_out_i_25_port, shifted_out_i_24_port, shifted_out_i_23_port, 
      shifted_out_i_22_port, shifted_out_i_21_port, shifted_out_i_20_port, 
      shifted_out_i_19_port, shifted_out_i_18_port, shifted_out_i_17_port, 
      shifted_out_i_16_port, shifted_out_i_15_port, shifted_out_i_14_port, 
      shifted_out_i_13_port, shifted_out_i_12_port, shifted_out_i_11_port, 
      shifted_out_i_10_port, shifted_out_i_9_port, shifted_out_i_8_port, 
      shifted_out_i_7_port, shifted_out_i_6_port, shifted_out_i_5_port, 
      shifted_out_i_4_port, shifted_out_i_3_port, shifted_out_i_2_port, 
      shifted_out_i_1_port, shifted_out_i_0_port : std_logic;

begin
   
   shifter_e : shifter_nbit32 port map( r1(31) => r1(31), r1(30) => r1(30), 
                           r1(29) => r1(29), r1(28) => r1(28), r1(27) => r1(27)
                           , r1(26) => r1(26), r1(25) => r1(25), r1(24) => 
                           r1(24), r1(23) => r1(23), r1(22) => r1(22), r1(21) 
                           => r1(21), r1(20) => r1(20), r1(19) => r1(19), 
                           r1(18) => r1(18), r1(17) => r1(17), r1(16) => r1(16)
                           , r1(15) => r1(15), r1(14) => r1(14), r1(13) => 
                           r1(13), r1(12) => r1(12), r1(11) => r1(11), r1(10) 
                           => r1(10), r1(9) => r1(9), r1(8) => r1(8), r1(7) => 
                           r1(7), r1(6) => r1(6), r1(5) => r1(5), r1(4) => 
                           r1(4), r1(3) => r1(3), r1(2) => r1(2), r1(1) => 
                           r1(1), r1(0) => r1(0), r2(31) => r2(31), r2(30) => 
                           r2(30), r2(29) => r2(29), r2(28) => r2(28), r2(27) 
                           => r2(27), r2(26) => r2(26), r2(25) => r2(25), 
                           r2(24) => r2(24), r2(23) => r2(23), r2(22) => r2(22)
                           , r2(21) => r2(21), r2(20) => r2(20), r2(19) => 
                           r2(19), r2(18) => r2(18), r2(17) => r2(17), r2(16) 
                           => r2(16), r2(15) => r2(15), r2(14) => r2(14), 
                           r2(13) => r2(13), r2(12) => r2(12), r2(11) => r2(11)
                           , r2(10) => r2(10), r2(9) => r2(9), r2(8) => r2(8), 
                           r2(7) => r2(7), r2(6) => r2(6), r2(5) => r2(5), 
                           r2(4) => r2(4), r2(3) => r2(3), r2(2) => r2(2), 
                           r2(1) => r2(1), r2(0) => r2(0), conf(1) => conf(1), 
                           conf(0) => conf(0), shifted_out(31) => 
                           shifted_out_i_31_port, shifted_out(30) => 
                           shifted_out_i_30_port, shifted_out(29) => 
                           shifted_out_i_29_port, shifted_out(28) => 
                           shifted_out_i_28_port, shifted_out(27) => 
                           shifted_out_i_27_port, shifted_out(26) => 
                           shifted_out_i_26_port, shifted_out(25) => 
                           shifted_out_i_25_port, shifted_out(24) => 
                           shifted_out_i_24_port, shifted_out(23) => 
                           shifted_out_i_23_port, shifted_out(22) => 
                           shifted_out_i_22_port, shifted_out(21) => 
                           shifted_out_i_21_port, shifted_out(20) => 
                           shifted_out_i_20_port, shifted_out(19) => 
                           shifted_out_i_19_port, shifted_out(18) => 
                           shifted_out_i_18_port, shifted_out(17) => 
                           shifted_out_i_17_port, shifted_out(16) => 
                           shifted_out_i_16_port, shifted_out(15) => 
                           shifted_out_i_15_port, shifted_out(14) => 
                           shifted_out_i_14_port, shifted_out(13) => 
                           shifted_out_i_13_port, shifted_out(12) => 
                           shifted_out_i_12_port, shifted_out(11) => 
                           shifted_out_i_11_port, shifted_out(10) => 
                           shifted_out_i_10_port, shifted_out(9) => 
                           shifted_out_i_9_port, shifted_out(8) => 
                           shifted_out_i_8_port, shifted_out(7) => 
                           shifted_out_i_7_port, shifted_out(6) => 
                           shifted_out_i_6_port, shifted_out(5) => 
                           shifted_out_i_5_port, shifted_out(4) => 
                           shifted_out_i_4_port, shifted_out(3) => 
                           shifted_out_i_3_port, shifted_out(2) => 
                           shifted_out_i_2_port, shifted_out(1) => 
                           shifted_out_i_1_port, shifted_out(0) => 
                           shifted_out_i_0_port);
   U2 : AND2_X1 port map( A1 => shifted_out_i_6_port, A2 => en_shifter, ZN => 
                           shifted_out(6));
   U3 : AND2_X1 port map( A1 => shifted_out_i_5_port, A2 => en_shifter, ZN => 
                           shifted_out(5));
   U4 : AND2_X1 port map( A1 => shifted_out_i_4_port, A2 => en_shifter, ZN => 
                           shifted_out(4));
   U5 : AND2_X1 port map( A1 => shifted_out_i_3_port, A2 => en_shifter, ZN => 
                           shifted_out(3));
   U6 : AND2_X1 port map( A1 => shifted_out_i_2_port, A2 => en_shifter, ZN => 
                           shifted_out(2));
   U7 : AND2_X1 port map( A1 => shifted_out_i_1_port, A2 => en_shifter, ZN => 
                           shifted_out(1));
   U8 : AND2_X1 port map( A1 => shifted_out_i_31_port, A2 => en_shifter, ZN => 
                           shifted_out(31));
   U9 : AND2_X1 port map( A1 => shifted_out_i_30_port, A2 => en_shifter, ZN => 
                           shifted_out(30));
   U10 : AND2_X1 port map( A1 => shifted_out_i_29_port, A2 => en_shifter, ZN =>
                           shifted_out(29));
   U11 : AND2_X1 port map( A1 => shifted_out_i_28_port, A2 => en_shifter, ZN =>
                           shifted_out(28));
   U12 : AND2_X1 port map( A1 => shifted_out_i_27_port, A2 => en_shifter, ZN =>
                           shifted_out(27));
   U13 : AND2_X1 port map( A1 => shifted_out_i_0_port, A2 => en_shifter, ZN => 
                           shifted_out(0));
   U14 : AND2_X1 port map( A1 => shifted_out_i_26_port, A2 => en_shifter, ZN =>
                           shifted_out(26));
   U15 : AND2_X1 port map( A1 => shifted_out_i_25_port, A2 => en_shifter, ZN =>
                           shifted_out(25));
   U16 : AND2_X1 port map( A1 => shifted_out_i_24_port, A2 => en_shifter, ZN =>
                           shifted_out(24));
   U17 : AND2_X1 port map( A1 => shifted_out_i_23_port, A2 => en_shifter, ZN =>
                           shifted_out(23));
   U18 : AND2_X1 port map( A1 => shifted_out_i_22_port, A2 => en_shifter, ZN =>
                           shifted_out(22));
   U19 : AND2_X1 port map( A1 => shifted_out_i_21_port, A2 => en_shifter, ZN =>
                           shifted_out(21));
   U20 : AND2_X1 port map( A1 => shifted_out_i_20_port, A2 => en_shifter, ZN =>
                           shifted_out(20));
   U21 : AND2_X1 port map( A1 => shifted_out_i_19_port, A2 => en_shifter, ZN =>
                           shifted_out(19));
   U22 : AND2_X1 port map( A1 => shifted_out_i_18_port, A2 => en_shifter, ZN =>
                           shifted_out(18));
   U23 : AND2_X1 port map( A1 => shifted_out_i_17_port, A2 => en_shifter, ZN =>
                           shifted_out(17));
   U24 : AND2_X1 port map( A1 => shifted_out_i_16_port, A2 => en_shifter, ZN =>
                           shifted_out(16));
   U25 : AND2_X1 port map( A1 => shifted_out_i_15_port, A2 => en_shifter, ZN =>
                           shifted_out(15));
   U26 : AND2_X1 port map( A1 => shifted_out_i_14_port, A2 => en_shifter, ZN =>
                           shifted_out(14));
   U27 : AND2_X1 port map( A1 => shifted_out_i_13_port, A2 => en_shifter, ZN =>
                           shifted_out(13));
   U28 : AND2_X1 port map( A1 => shifted_out_i_12_port, A2 => en_shifter, ZN =>
                           shifted_out(12));
   U29 : AND2_X1 port map( A1 => shifted_out_i_11_port, A2 => en_shifter, ZN =>
                           shifted_out(11));
   U30 : AND2_X1 port map( A1 => shifted_out_i_10_port, A2 => en_shifter, ZN =>
                           shifted_out(10));
   U31 : AND2_X1 port map( A1 => shifted_out_i_9_port, A2 => en_shifter, ZN => 
                           shifted_out(9));
   U32 : AND2_X1 port map( A1 => shifted_out_i_8_port, A2 => en_shifter, ZN => 
                           shifted_out(8));
   U33 : AND2_X1 port map( A1 => shifted_out_i_7_port, A2 => en_shifter, ZN => 
                           shifted_out(7));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity zero_comparator_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  en : in std_logic;  cond : 
         in std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
         0));

end zero_comparator_N32;

architecture SYN_Behavioral of zero_comparator_N32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component zero_comparator_N32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal O_31_port, N68, N70, N72, n10, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n_1426, n_1427, 
      n_1428 : std_logic;

begin
   O <= ( O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, 
      O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, 
      O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, 
      O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, 
      O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, O_31_port, 
      O_31_port, O_31_port );
   
   n10 <= '0';
   r70 : zero_comparator_N32_DW01_cmp6_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), TC => n10, LT => N72, GT => 
                           N70, EQ => n_1426, LE => n_1427, GE => n_1428, NE =>
                           N68);
   U3 : AND2_X1 port map( A1 => n1, A2 => en, ZN => O_31_port);
   U4 : MUX2_X1 port map( A => n2, B => n3, S => cond(2), Z => n1);
   U5 : MUX2_X1 port map( A => n4, B => n5, S => cond(1), Z => n3);
   U6 : NOR2_X1 port map( A1 => cond(0), A2 => n6, ZN => n5);
   U7 : XOR2_X1 port map( A => N70, B => cond(0), Z => n4);
   U8 : MUX2_X1 port map( A => n7, B => n8, S => cond(1), Z => n2);
   U9 : MUX2_X1 port map( A => N68, B => n6, S => cond(0), Z => n8);
   U10 : INV_X1 port map( A => N72, ZN => n6);
   U11 : MUX2_X1 port map( A => n9, B => n11, S => cond(0), Z => n7);
   U12 : INV_X1 port map( A => N68, ZN => n11);
   U13 : NOR2_X1 port map( A1 => n12, A2 => n13, ZN => n9);
   U14 : NAND4_X1 port map( A1 => n14, A2 => n15, A3 => n16, A4 => n17, ZN => 
                           n13);
   U15 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n17);
   U16 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), 
                           ZN => n16);
   U17 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n15);
   U18 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), 
                           ZN => n14);
   U19 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n12);
   U20 : NOR4_X1 port map( A1 => A(9), A2 => A(8), A3 => A(7), A4 => A(6), ZN 
                           => n21);
   U21 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n20);
   U22 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), 
                           ZN => n19);
   U23 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n18);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity mul_wrapper_NBIT32_N16_M16 is

   port( a, b : in std_logic_vector (31 downto 0);  en : in std_logic;  mul : 
         out std_logic_vector (31 downto 0));

end mul_wrapper_NBIT32_N16_M16;

architecture SYN_specification of mul_wrapper_NBIT32_N16_M16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component boothmul_NBIT32_N16_M16
      port( a, b : in std_logic_vector (15 downto 0);  mul : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal mul_out_31_port, mul_out_30_port, mul_out_29_port, mul_out_28_port, 
      mul_out_27_port, mul_out_26_port, mul_out_25_port, mul_out_24_port, 
      mul_out_23_port, mul_out_22_port, mul_out_21_port, mul_out_20_port, 
      mul_out_19_port, mul_out_18_port, mul_out_17_port, mul_out_16_port, 
      mul_out_15_port, mul_out_14_port, mul_out_13_port, mul_out_12_port, 
      mul_out_11_port, mul_out_10_port, mul_out_9_port, mul_out_8_port, 
      mul_out_7_port, mul_out_6_port, mul_out_5_port, mul_out_4_port, 
      mul_out_3_port, mul_out_2_port, mul_out_1_port, mul_out_0_port : 
      std_logic;

begin
   
   mult : boothmul_NBIT32_N16_M16 port map( a(15) => a(15), a(14) => a(14), 
                           a(13) => a(13), a(12) => a(12), a(11) => a(11), 
                           a(10) => a(10), a(9) => a(9), a(8) => a(8), a(7) => 
                           a(7), a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3)
                           => a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), mul(31) => 
                           mul_out_31_port, mul(30) => mul_out_30_port, mul(29)
                           => mul_out_29_port, mul(28) => mul_out_28_port, 
                           mul(27) => mul_out_27_port, mul(26) => 
                           mul_out_26_port, mul(25) => mul_out_25_port, mul(24)
                           => mul_out_24_port, mul(23) => mul_out_23_port, 
                           mul(22) => mul_out_22_port, mul(21) => 
                           mul_out_21_port, mul(20) => mul_out_20_port, mul(19)
                           => mul_out_19_port, mul(18) => mul_out_18_port, 
                           mul(17) => mul_out_17_port, mul(16) => 
                           mul_out_16_port, mul(15) => mul_out_15_port, mul(14)
                           => mul_out_14_port, mul(13) => mul_out_13_port, 
                           mul(12) => mul_out_12_port, mul(11) => 
                           mul_out_11_port, mul(10) => mul_out_10_port, mul(9) 
                           => mul_out_9_port, mul(8) => mul_out_8_port, mul(7) 
                           => mul_out_7_port, mul(6) => mul_out_6_port, mul(5) 
                           => mul_out_5_port, mul(4) => mul_out_4_port, mul(3) 
                           => mul_out_3_port, mul(2) => mul_out_2_port, mul(1) 
                           => mul_out_1_port, mul(0) => mul_out_0_port);
   U2 : AND2_X1 port map( A1 => mul_out_9_port, A2 => en, ZN => mul(9));
   U3 : AND2_X1 port map( A1 => mul_out_8_port, A2 => en, ZN => mul(8));
   U4 : AND2_X1 port map( A1 => mul_out_7_port, A2 => en, ZN => mul(7));
   U5 : AND2_X1 port map( A1 => mul_out_6_port, A2 => en, ZN => mul(6));
   U6 : AND2_X1 port map( A1 => mul_out_5_port, A2 => en, ZN => mul(5));
   U7 : AND2_X1 port map( A1 => mul_out_4_port, A2 => en, ZN => mul(4));
   U8 : AND2_X1 port map( A1 => mul_out_3_port, A2 => en, ZN => mul(3));
   U9 : AND2_X1 port map( A1 => mul_out_31_port, A2 => en, ZN => mul(31));
   U10 : AND2_X1 port map( A1 => mul_out_30_port, A2 => en, ZN => mul(30));
   U11 : AND2_X1 port map( A1 => mul_out_2_port, A2 => en, ZN => mul(2));
   U12 : AND2_X1 port map( A1 => mul_out_29_port, A2 => en, ZN => mul(29));
   U13 : AND2_X1 port map( A1 => mul_out_28_port, A2 => en, ZN => mul(28));
   U14 : AND2_X1 port map( A1 => mul_out_27_port, A2 => en, ZN => mul(27));
   U15 : AND2_X1 port map( A1 => mul_out_26_port, A2 => en, ZN => mul(26));
   U16 : AND2_X1 port map( A1 => mul_out_25_port, A2 => en, ZN => mul(25));
   U17 : AND2_X1 port map( A1 => mul_out_24_port, A2 => en, ZN => mul(24));
   U18 : AND2_X1 port map( A1 => mul_out_23_port, A2 => en, ZN => mul(23));
   U19 : AND2_X1 port map( A1 => mul_out_22_port, A2 => en, ZN => mul(22));
   U20 : AND2_X1 port map( A1 => mul_out_21_port, A2 => en, ZN => mul(21));
   U21 : AND2_X1 port map( A1 => mul_out_20_port, A2 => en, ZN => mul(20));
   U22 : AND2_X1 port map( A1 => mul_out_1_port, A2 => en, ZN => mul(1));
   U23 : AND2_X1 port map( A1 => mul_out_19_port, A2 => en, ZN => mul(19));
   U24 : AND2_X1 port map( A1 => mul_out_18_port, A2 => en, ZN => mul(18));
   U25 : AND2_X1 port map( A1 => mul_out_17_port, A2 => en, ZN => mul(17));
   U26 : AND2_X1 port map( A1 => mul_out_16_port, A2 => en, ZN => mul(16));
   U27 : AND2_X1 port map( A1 => mul_out_15_port, A2 => en, ZN => mul(15));
   U28 : AND2_X1 port map( A1 => mul_out_14_port, A2 => en, ZN => mul(14));
   U29 : AND2_X1 port map( A1 => mul_out_13_port, A2 => en, ZN => mul(13));
   U30 : AND2_X1 port map( A1 => mul_out_12_port, A2 => en, ZN => mul(12));
   U31 : AND2_X1 port map( A1 => mul_out_11_port, A2 => en, ZN => mul(11));
   U32 : AND2_X1 port map( A1 => mul_out_10_port, A2 => en, ZN => mul(10));
   U33 : AND2_X1 port map( A1 => mul_out_0_port, A2 => en, ZN => mul(0));

end SYN_specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity adder_wrapper_nbit32 is

   port( op1, op2 : in std_logic_vector (31 downto 0);  CarryIn : in std_logic;
         sum : out std_logic_vector (31 downto 0);  CarryOut, overflow : out 
         std_logic;  en_adder : in std_logic);

end adder_wrapper_nbit32;

architecture SYN_Behavioral of adder_wrapper_nbit32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sparse_tree_adder_n_bit32
      port( operand_1, operand_2 : in std_logic_vector (31 downto 0);  carry_in
            : in std_logic;  sum : out std_logic_vector (31 downto 0);  
            carry_out, overflow : out std_logic);
   end component;
   
   component MUX21_N32_1
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal op2_mux_31_port, op2_mux_30_port, op2_mux_29_port, op2_mux_28_port, 
      op2_mux_27_port, op2_mux_26_port, op2_mux_25_port, op2_mux_24_port, 
      op2_mux_23_port, op2_mux_22_port, op2_mux_21_port, op2_mux_20_port, 
      op2_mux_19_port, op2_mux_18_port, op2_mux_17_port, op2_mux_16_port, 
      op2_mux_15_port, op2_mux_14_port, op2_mux_13_port, op2_mux_12_port, 
      op2_mux_11_port, op2_mux_10_port, op2_mux_9_port, op2_mux_8_port, 
      op2_mux_7_port, op2_mux_6_port, op2_mux_5_port, op2_mux_4_port, 
      op2_mux_3_port, op2_mux_2_port, op2_mux_1_port, op2_mux_0_port, 
      sum_out_31_port, sum_out_30_port, sum_out_29_port, sum_out_28_port, 
      sum_out_27_port, sum_out_26_port, sum_out_25_port, sum_out_24_port, 
      sum_out_23_port, sum_out_22_port, sum_out_21_port, sum_out_20_port, 
      sum_out_19_port, sum_out_18_port, sum_out_17_port, sum_out_16_port, 
      sum_out_15_port, sum_out_14_port, sum_out_13_port, sum_out_12_port, 
      sum_out_11_port, sum_out_10_port, sum_out_9_port, sum_out_8_port, 
      sum_out_7_port, sum_out_6_port, sum_out_5_port, sum_out_4_port, 
      sum_out_3_port, sum_out_2_port, sum_out_1_port, sum_out_0_port, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32 : 
      std_logic;

begin
   
   mux_operand2 : MUX21_N32_1 port map( a(31) => op2(31), a(30) => op2(30), 
                           a(29) => op2(29), a(28) => op2(28), a(27) => op2(27)
                           , a(26) => op2(26), a(25) => op2(25), a(24) => 
                           op2(24), a(23) => op2(23), a(22) => op2(22), a(21) 
                           => op2(21), a(20) => op2(20), a(19) => op2(19), 
                           a(18) => op2(18), a(17) => op2(17), a(16) => op2(16)
                           , a(15) => op2(15), a(14) => op2(14), a(13) => 
                           op2(13), a(12) => op2(12), a(11) => op2(11), a(10) 
                           => op2(10), a(9) => op2(9), a(8) => op2(8), a(7) => 
                           op2(7), a(6) => op2(6), a(5) => op2(5), a(4) => 
                           op2(4), a(3) => op2(3), a(2) => op2(2), a(1) => 
                           op2(1), a(0) => op2(0), b(31) => n1, b(30) => n2, 
                           b(29) => n3, b(28) => n4, b(27) => n5, b(26) => n6, 
                           b(25) => n7, b(24) => n8, b(23) => n9, b(22) => n10,
                           b(21) => n11, b(20) => n12, b(19) => n13, b(18) => 
                           n14, b(17) => n15, b(16) => n16, b(15) => n17, b(14)
                           => n18, b(13) => n19, b(12) => n20, b(11) => n21, 
                           b(10) => n22, b(9) => n23, b(8) => n24, b(7) => n25,
                           b(6) => n26, b(5) => n27, b(4) => n28, b(3) => n29, 
                           b(2) => n30, b(1) => n31, b(0) => n32, sel => 
                           CarryIn, y(31) => op2_mux_31_port, y(30) => 
                           op2_mux_30_port, y(29) => op2_mux_29_port, y(28) => 
                           op2_mux_28_port, y(27) => op2_mux_27_port, y(26) => 
                           op2_mux_26_port, y(25) => op2_mux_25_port, y(24) => 
                           op2_mux_24_port, y(23) => op2_mux_23_port, y(22) => 
                           op2_mux_22_port, y(21) => op2_mux_21_port, y(20) => 
                           op2_mux_20_port, y(19) => op2_mux_19_port, y(18) => 
                           op2_mux_18_port, y(17) => op2_mux_17_port, y(16) => 
                           op2_mux_16_port, y(15) => op2_mux_15_port, y(14) => 
                           op2_mux_14_port, y(13) => op2_mux_13_port, y(12) => 
                           op2_mux_12_port, y(11) => op2_mux_11_port, y(10) => 
                           op2_mux_10_port, y(9) => op2_mux_9_port, y(8) => 
                           op2_mux_8_port, y(7) => op2_mux_7_port, y(6) => 
                           op2_mux_6_port, y(5) => op2_mux_5_port, y(4) => 
                           op2_mux_4_port, y(3) => op2_mux_3_port, y(2) => 
                           op2_mux_2_port, y(1) => op2_mux_1_port, y(0) => 
                           op2_mux_0_port);
   sparse_adder : sparse_tree_adder_n_bit32 port map( operand_1(31) => op1(31),
                           operand_1(30) => op1(30), operand_1(29) => op1(29), 
                           operand_1(28) => op1(28), operand_1(27) => op1(27), 
                           operand_1(26) => op1(26), operand_1(25) => op1(25), 
                           operand_1(24) => op1(24), operand_1(23) => op1(23), 
                           operand_1(22) => op1(22), operand_1(21) => op1(21), 
                           operand_1(20) => op1(20), operand_1(19) => op1(19), 
                           operand_1(18) => op1(18), operand_1(17) => op1(17), 
                           operand_1(16) => op1(16), operand_1(15) => op1(15), 
                           operand_1(14) => op1(14), operand_1(13) => op1(13), 
                           operand_1(12) => op1(12), operand_1(11) => op1(11), 
                           operand_1(10) => op1(10), operand_1(9) => op1(9), 
                           operand_1(8) => op1(8), operand_1(7) => op1(7), 
                           operand_1(6) => op1(6), operand_1(5) => op1(5), 
                           operand_1(4) => op1(4), operand_1(3) => op1(3), 
                           operand_1(2) => op1(2), operand_1(1) => op1(1), 
                           operand_1(0) => op1(0), operand_2(31) => 
                           op2_mux_31_port, operand_2(30) => op2_mux_30_port, 
                           operand_2(29) => op2_mux_29_port, operand_2(28) => 
                           op2_mux_28_port, operand_2(27) => op2_mux_27_port, 
                           operand_2(26) => op2_mux_26_port, operand_2(25) => 
                           op2_mux_25_port, operand_2(24) => op2_mux_24_port, 
                           operand_2(23) => op2_mux_23_port, operand_2(22) => 
                           op2_mux_22_port, operand_2(21) => op2_mux_21_port, 
                           operand_2(20) => op2_mux_20_port, operand_2(19) => 
                           op2_mux_19_port, operand_2(18) => op2_mux_18_port, 
                           operand_2(17) => op2_mux_17_port, operand_2(16) => 
                           op2_mux_16_port, operand_2(15) => op2_mux_15_port, 
                           operand_2(14) => op2_mux_14_port, operand_2(13) => 
                           op2_mux_13_port, operand_2(12) => op2_mux_12_port, 
                           operand_2(11) => op2_mux_11_port, operand_2(10) => 
                           op2_mux_10_port, operand_2(9) => op2_mux_9_port, 
                           operand_2(8) => op2_mux_8_port, operand_2(7) => 
                           op2_mux_7_port, operand_2(6) => op2_mux_6_port, 
                           operand_2(5) => op2_mux_5_port, operand_2(4) => 
                           op2_mux_4_port, operand_2(3) => op2_mux_3_port, 
                           operand_2(2) => op2_mux_2_port, operand_2(1) => 
                           op2_mux_1_port, operand_2(0) => op2_mux_0_port, 
                           carry_in => CarryIn, sum(31) => sum_out_31_port, 
                           sum(30) => sum_out_30_port, sum(29) => 
                           sum_out_29_port, sum(28) => sum_out_28_port, sum(27)
                           => sum_out_27_port, sum(26) => sum_out_26_port, 
                           sum(25) => sum_out_25_port, sum(24) => 
                           sum_out_24_port, sum(23) => sum_out_23_port, sum(22)
                           => sum_out_22_port, sum(21) => sum_out_21_port, 
                           sum(20) => sum_out_20_port, sum(19) => 
                           sum_out_19_port, sum(18) => sum_out_18_port, sum(17)
                           => sum_out_17_port, sum(16) => sum_out_16_port, 
                           sum(15) => sum_out_15_port, sum(14) => 
                           sum_out_14_port, sum(13) => sum_out_13_port, sum(12)
                           => sum_out_12_port, sum(11) => sum_out_11_port, 
                           sum(10) => sum_out_10_port, sum(9) => sum_out_9_port
                           , sum(8) => sum_out_8_port, sum(7) => sum_out_7_port
                           , sum(6) => sum_out_6_port, sum(5) => sum_out_5_port
                           , sum(4) => sum_out_4_port, sum(3) => sum_out_3_port
                           , sum(2) => sum_out_2_port, sum(1) => sum_out_1_port
                           , sum(0) => sum_out_0_port, carry_out => CarryOut, 
                           overflow => overflow);
   U2 : AND2_X1 port map( A1 => sum_out_9_port, A2 => en_adder, ZN => sum(9));
   U3 : AND2_X1 port map( A1 => sum_out_8_port, A2 => en_adder, ZN => sum(8));
   U4 : AND2_X1 port map( A1 => sum_out_7_port, A2 => en_adder, ZN => sum(7));
   U5 : AND2_X1 port map( A1 => sum_out_6_port, A2 => en_adder, ZN => sum(6));
   U6 : AND2_X1 port map( A1 => sum_out_5_port, A2 => en_adder, ZN => sum(5));
   U7 : AND2_X1 port map( A1 => sum_out_4_port, A2 => en_adder, ZN => sum(4));
   U8 : AND2_X1 port map( A1 => sum_out_3_port, A2 => en_adder, ZN => sum(3));
   U9 : AND2_X1 port map( A1 => sum_out_31_port, A2 => en_adder, ZN => sum(31))
                           ;
   U10 : AND2_X1 port map( A1 => sum_out_30_port, A2 => en_adder, ZN => sum(30)
                           );
   U11 : AND2_X1 port map( A1 => sum_out_2_port, A2 => en_adder, ZN => sum(2));
   U12 : AND2_X1 port map( A1 => sum_out_29_port, A2 => en_adder, ZN => sum(29)
                           );
   U13 : AND2_X1 port map( A1 => sum_out_28_port, A2 => en_adder, ZN => sum(28)
                           );
   U14 : AND2_X1 port map( A1 => sum_out_27_port, A2 => en_adder, ZN => sum(27)
                           );
   U15 : AND2_X1 port map( A1 => sum_out_26_port, A2 => en_adder, ZN => sum(26)
                           );
   U16 : AND2_X1 port map( A1 => sum_out_25_port, A2 => en_adder, ZN => sum(25)
                           );
   U17 : AND2_X1 port map( A1 => sum_out_24_port, A2 => en_adder, ZN => sum(24)
                           );
   U18 : AND2_X1 port map( A1 => sum_out_23_port, A2 => en_adder, ZN => sum(23)
                           );
   U19 : AND2_X1 port map( A1 => sum_out_22_port, A2 => en_adder, ZN => sum(22)
                           );
   U20 : AND2_X1 port map( A1 => sum_out_21_port, A2 => en_adder, ZN => sum(21)
                           );
   U21 : AND2_X1 port map( A1 => sum_out_20_port, A2 => en_adder, ZN => sum(20)
                           );
   U22 : AND2_X1 port map( A1 => sum_out_1_port, A2 => en_adder, ZN => sum(1));
   U23 : AND2_X1 port map( A1 => sum_out_19_port, A2 => en_adder, ZN => sum(19)
                           );
   U24 : AND2_X1 port map( A1 => sum_out_18_port, A2 => en_adder, ZN => sum(18)
                           );
   U25 : AND2_X1 port map( A1 => sum_out_17_port, A2 => en_adder, ZN => sum(17)
                           );
   U26 : AND2_X1 port map( A1 => sum_out_16_port, A2 => en_adder, ZN => sum(16)
                           );
   U27 : AND2_X1 port map( A1 => sum_out_15_port, A2 => en_adder, ZN => sum(15)
                           );
   U28 : AND2_X1 port map( A1 => sum_out_14_port, A2 => en_adder, ZN => sum(14)
                           );
   U29 : AND2_X1 port map( A1 => sum_out_13_port, A2 => en_adder, ZN => sum(13)
                           );
   U30 : AND2_X1 port map( A1 => sum_out_12_port, A2 => en_adder, ZN => sum(12)
                           );
   U31 : AND2_X1 port map( A1 => sum_out_11_port, A2 => en_adder, ZN => sum(11)
                           );
   U32 : AND2_X1 port map( A1 => sum_out_10_port, A2 => en_adder, ZN => sum(10)
                           );
   U33 : AND2_X1 port map( A1 => sum_out_0_port, A2 => en_adder, ZN => sum(0));
   U34 : INV_X1 port map( A => op2(31), ZN => n1);
   U35 : INV_X1 port map( A => op2(30), ZN => n2);
   U36 : INV_X1 port map( A => op2(29), ZN => n3);
   U37 : INV_X1 port map( A => op2(28), ZN => n4);
   U38 : INV_X1 port map( A => op2(27), ZN => n5);
   U39 : INV_X1 port map( A => op2(26), ZN => n6);
   U40 : INV_X1 port map( A => op2(25), ZN => n7);
   U41 : INV_X1 port map( A => op2(24), ZN => n8);
   U42 : INV_X1 port map( A => op2(23), ZN => n9);
   U43 : INV_X1 port map( A => op2(22), ZN => n10);
   U44 : INV_X1 port map( A => op2(21), ZN => n11);
   U45 : INV_X1 port map( A => op2(20), ZN => n12);
   U46 : INV_X1 port map( A => op2(19), ZN => n13);
   U47 : INV_X1 port map( A => op2(18), ZN => n14);
   U48 : INV_X1 port map( A => op2(17), ZN => n15);
   U49 : INV_X1 port map( A => op2(16), ZN => n16);
   U50 : INV_X1 port map( A => op2(15), ZN => n17);
   U51 : INV_X1 port map( A => op2(14), ZN => n18);
   U52 : INV_X1 port map( A => op2(13), ZN => n19);
   U53 : INV_X1 port map( A => op2(12), ZN => n20);
   U54 : INV_X1 port map( A => op2(11), ZN => n21);
   U55 : INV_X1 port map( A => op2(10), ZN => n22);
   U56 : INV_X1 port map( A => op2(9), ZN => n23);
   U57 : INV_X1 port map( A => op2(8), ZN => n24);
   U58 : INV_X1 port map( A => op2(7), ZN => n25);
   U59 : INV_X1 port map( A => op2(6), ZN => n26);
   U60 : INV_X1 port map( A => op2(5), ZN => n27);
   U61 : INV_X1 port map( A => op2(4), ZN => n28);
   U62 : INV_X1 port map( A => op2(3), ZN => n29);
   U63 : INV_X1 port map( A => op2(2), ZN => n30);
   U64 : INV_X1 port map( A => op2(1), ZN => n31);
   U65 : INV_X1 port map( A => op2(0), ZN => n32);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity logic_op_unit_Nbit32 is

   port( op1, op2 : in std_logic_vector (31 downto 0);  en_logic, s3, s2, s1, 
         s0 : in std_logic;  logic_out : out std_logic_vector (31 downto 0));

end logic_op_unit_Nbit32;

architecture SYN_logic_op_unit_arc of logic_op_unit_Nbit32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => n1, B => n2, S => op2(9), Z => logic_out(9));
   U2 : MUX2_X1 port map( A => s1, B => s3, S => op1(9), Z => n2);
   U3 : MUX2_X1 port map( A => s0, B => s2, S => op1(9), Z => n1);
   U4 : MUX2_X1 port map( A => n3, B => n4, S => op2(8), Z => logic_out(8));
   U5 : MUX2_X1 port map( A => s1, B => s3, S => op1(8), Z => n4);
   U6 : MUX2_X1 port map( A => s0, B => s2, S => op1(8), Z => n3);
   U7 : MUX2_X1 port map( A => n5, B => n6, S => op2(7), Z => logic_out(7));
   U8 : MUX2_X1 port map( A => s1, B => s3, S => op1(7), Z => n6);
   U9 : MUX2_X1 port map( A => s0, B => s2, S => op1(7), Z => n5);
   U10 : MUX2_X1 port map( A => n7, B => n8, S => op2(6), Z => logic_out(6));
   U11 : MUX2_X1 port map( A => s1, B => s3, S => op1(6), Z => n8);
   U12 : MUX2_X1 port map( A => s0, B => s2, S => op1(6), Z => n7);
   U13 : MUX2_X1 port map( A => n9, B => n10, S => op2(5), Z => logic_out(5));
   U14 : MUX2_X1 port map( A => s1, B => s3, S => op1(5), Z => n10);
   U15 : MUX2_X1 port map( A => s0, B => s2, S => op1(5), Z => n9);
   U16 : MUX2_X1 port map( A => n11, B => n12, S => op2(4), Z => logic_out(4));
   U17 : MUX2_X1 port map( A => s1, B => s3, S => op1(4), Z => n12);
   U18 : MUX2_X1 port map( A => s0, B => s2, S => op1(4), Z => n11);
   U19 : MUX2_X1 port map( A => n13, B => n14, S => op2(3), Z => logic_out(3));
   U20 : MUX2_X1 port map( A => s1, B => s3, S => op1(3), Z => n14);
   U21 : MUX2_X1 port map( A => s0, B => s2, S => op1(3), Z => n13);
   U22 : MUX2_X1 port map( A => n15, B => n16, S => op2(31), Z => logic_out(31)
                           );
   U23 : MUX2_X1 port map( A => s1, B => s3, S => op1(31), Z => n16);
   U24 : MUX2_X1 port map( A => s0, B => s2, S => op1(31), Z => n15);
   U25 : MUX2_X1 port map( A => n17, B => n18, S => op2(30), Z => logic_out(30)
                           );
   U26 : MUX2_X1 port map( A => s1, B => s3, S => op1(30), Z => n18);
   U27 : MUX2_X1 port map( A => s0, B => s2, S => op1(30), Z => n17);
   U28 : MUX2_X1 port map( A => n19, B => n20, S => op2(2), Z => logic_out(2));
   U29 : MUX2_X1 port map( A => s1, B => s3, S => op1(2), Z => n20);
   U30 : MUX2_X1 port map( A => s0, B => s2, S => op1(2), Z => n19);
   U31 : MUX2_X1 port map( A => n21, B => n22, S => op2(29), Z => logic_out(29)
                           );
   U32 : MUX2_X1 port map( A => s1, B => s3, S => op1(29), Z => n22);
   U33 : MUX2_X1 port map( A => s0, B => s2, S => op1(29), Z => n21);
   U34 : MUX2_X1 port map( A => n23, B => n24, S => op2(28), Z => logic_out(28)
                           );
   U35 : MUX2_X1 port map( A => s1, B => s3, S => op1(28), Z => n24);
   U36 : MUX2_X1 port map( A => s0, B => s2, S => op1(28), Z => n23);
   U37 : MUX2_X1 port map( A => n25, B => n26, S => op2(27), Z => logic_out(27)
                           );
   U38 : MUX2_X1 port map( A => s1, B => s3, S => op1(27), Z => n26);
   U39 : MUX2_X1 port map( A => s0, B => s2, S => op1(27), Z => n25);
   U40 : MUX2_X1 port map( A => n27, B => n28, S => op2(26), Z => logic_out(26)
                           );
   U41 : MUX2_X1 port map( A => s1, B => s3, S => op1(26), Z => n28);
   U42 : MUX2_X1 port map( A => s0, B => s2, S => op1(26), Z => n27);
   U43 : MUX2_X1 port map( A => n29, B => n30, S => op2(25), Z => logic_out(25)
                           );
   U44 : MUX2_X1 port map( A => s1, B => s3, S => op1(25), Z => n30);
   U45 : MUX2_X1 port map( A => s0, B => s2, S => op1(25), Z => n29);
   U46 : MUX2_X1 port map( A => n31, B => n32, S => op2(24), Z => logic_out(24)
                           );
   U47 : MUX2_X1 port map( A => s1, B => s3, S => op1(24), Z => n32);
   U48 : MUX2_X1 port map( A => s0, B => s2, S => op1(24), Z => n31);
   U49 : MUX2_X1 port map( A => n33, B => n34, S => op2(23), Z => logic_out(23)
                           );
   U50 : MUX2_X1 port map( A => s1, B => s3, S => op1(23), Z => n34);
   U51 : MUX2_X1 port map( A => s0, B => s2, S => op1(23), Z => n33);
   U52 : MUX2_X1 port map( A => n35, B => n36, S => op2(22), Z => logic_out(22)
                           );
   U53 : MUX2_X1 port map( A => s1, B => s3, S => op1(22), Z => n36);
   U54 : MUX2_X1 port map( A => s0, B => s2, S => op1(22), Z => n35);
   U55 : MUX2_X1 port map( A => n37, B => n38, S => op2(21), Z => logic_out(21)
                           );
   U56 : MUX2_X1 port map( A => s1, B => s3, S => op1(21), Z => n38);
   U57 : MUX2_X1 port map( A => s0, B => s2, S => op1(21), Z => n37);
   U58 : MUX2_X1 port map( A => n39, B => n40, S => op2(20), Z => logic_out(20)
                           );
   U59 : MUX2_X1 port map( A => s1, B => s3, S => op1(20), Z => n40);
   U60 : MUX2_X1 port map( A => s0, B => s2, S => op1(20), Z => n39);
   U61 : MUX2_X1 port map( A => n41, B => n42, S => op2(1), Z => logic_out(1));
   U62 : MUX2_X1 port map( A => s1, B => s3, S => op1(1), Z => n42);
   U63 : MUX2_X1 port map( A => s0, B => s2, S => op1(1), Z => n41);
   U64 : MUX2_X1 port map( A => n43, B => n44, S => op2(19), Z => logic_out(19)
                           );
   U65 : MUX2_X1 port map( A => s1, B => s3, S => op1(19), Z => n44);
   U66 : MUX2_X1 port map( A => s0, B => s2, S => op1(19), Z => n43);
   U67 : MUX2_X1 port map( A => n45, B => n46, S => op2(18), Z => logic_out(18)
                           );
   U68 : MUX2_X1 port map( A => s1, B => s3, S => op1(18), Z => n46);
   U69 : MUX2_X1 port map( A => s0, B => s2, S => op1(18), Z => n45);
   U70 : MUX2_X1 port map( A => n47, B => n48, S => op2(17), Z => logic_out(17)
                           );
   U71 : MUX2_X1 port map( A => s1, B => s3, S => op1(17), Z => n48);
   U72 : MUX2_X1 port map( A => s0, B => s2, S => op1(17), Z => n47);
   U73 : MUX2_X1 port map( A => n49, B => n50, S => op2(16), Z => logic_out(16)
                           );
   U74 : MUX2_X1 port map( A => s1, B => s3, S => op1(16), Z => n50);
   U75 : MUX2_X1 port map( A => s0, B => s2, S => op1(16), Z => n49);
   U76 : MUX2_X1 port map( A => n51, B => n52, S => op2(15), Z => logic_out(15)
                           );
   U77 : MUX2_X1 port map( A => s1, B => s3, S => op1(15), Z => n52);
   U78 : MUX2_X1 port map( A => s0, B => s2, S => op1(15), Z => n51);
   U79 : MUX2_X1 port map( A => n53, B => n54, S => op2(14), Z => logic_out(14)
                           );
   U80 : MUX2_X1 port map( A => s1, B => s3, S => op1(14), Z => n54);
   U81 : MUX2_X1 port map( A => s0, B => s2, S => op1(14), Z => n53);
   U82 : MUX2_X1 port map( A => n55, B => n56, S => op2(13), Z => logic_out(13)
                           );
   U83 : MUX2_X1 port map( A => s1, B => s3, S => op1(13), Z => n56);
   U84 : MUX2_X1 port map( A => s0, B => s2, S => op1(13), Z => n55);
   U85 : MUX2_X1 port map( A => n57, B => n58, S => op2(12), Z => logic_out(12)
                           );
   U86 : MUX2_X1 port map( A => s1, B => s3, S => op1(12), Z => n58);
   U87 : MUX2_X1 port map( A => s0, B => s2, S => op1(12), Z => n57);
   U88 : MUX2_X1 port map( A => n59, B => n60, S => op2(11), Z => logic_out(11)
                           );
   U89 : MUX2_X1 port map( A => s1, B => s3, S => op1(11), Z => n60);
   U90 : MUX2_X1 port map( A => s0, B => s2, S => op1(11), Z => n59);
   U91 : MUX2_X1 port map( A => n61, B => n62, S => op2(10), Z => logic_out(10)
                           );
   U92 : MUX2_X1 port map( A => s1, B => s3, S => op1(10), Z => n62);
   U93 : MUX2_X1 port map( A => s0, B => s2, S => op1(10), Z => n61);
   U94 : MUX2_X1 port map( A => n63, B => n64, S => op2(0), Z => logic_out(0));
   U95 : MUX2_X1 port map( A => s1, B => s3, S => op1(0), Z => n64);
   U96 : MUX2_X1 port map( A => s0, B => s2, S => op1(0), Z => n63);

end SYN_logic_op_unit_arc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ALU_decoder is

   port( s5, s4, s3, s2, s1, s0, en_ALU : in std_logic;  en_mult, en_comp, 
         en_Shift, en_Adder, en_Logic : out std_logic);

end ALU_decoder;

architecture SYN_ALU_decoder_beh of ALU_decoder is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n10 : std_logic;

begin
   
   U2 : OR3_X1 port map( A1 => n7, A2 => s5, A3 => n10, ZN => n1);
   U3 : OR2_X1 port map( A1 => s4, A2 => n8, ZN => n2);
   U4 : OR3_X1 port map( A1 => n7, A2 => n8, A3 => n9, ZN => n3);
   U5 : INV_X1 port map( A => n2, ZN => en_Shift);
   U6 : INV_X1 port map( A => n1, ZN => en_Adder);
   U7 : INV_X4 port map( A => n3, ZN => en_mult);
   U8 : INV_X1 port map( A => s3, ZN => n9);
   U9 : NOR3_X1 port map( A1 => n7, A2 => s3, A3 => n8, ZN => en_comp);
   U10 : NAND2_X1 port map( A1 => s5, A2 => en_ALU, ZN => n8);
   U11 : NOR3_X1 port map( A1 => n10, A2 => s5, A3 => s4, ZN => en_Logic);
   U12 : INV_X1 port map( A => en_ALU, ZN => n10);
   U13 : INV_X1 port map( A => s4, ZN => n7);

end SYN_ALU_decoder_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity ALU_NBIT32 is

   port( en_alu : in std_logic;  op1, op2 : in std_logic_vector (31 downto 0); 
         sel : in std_logic_vector (5 downto 0);  result : out std_logic_vector
         (31 downto 0);  CarryOut, overflow : out std_logic);

end ALU_NBIT32;

architecture SYN_Specification of ALU_NBIT32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shifter_wrapper_nbit32
      port( r1, r2 : in std_logic_vector (31 downto 0);  conf : in 
            std_logic_vector (1 downto 0);  en_shifter : in std_logic;  
            shifted_out : out std_logic_vector (31 downto 0));
   end component;
   
   component zero_comparator_N32
      port( A, B : in std_logic_vector (31 downto 0);  en : in std_logic;  cond
            : in std_logic_vector (2 downto 0);  O : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mul_wrapper_NBIT32_N16_M16
      port( a, b : in std_logic_vector (31 downto 0);  en : in std_logic;  mul 
            : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_wrapper_nbit32
      port( op1, op2 : in std_logic_vector (31 downto 0);  CarryIn : in 
            std_logic;  sum : out std_logic_vector (31 downto 0);  CarryOut, 
            overflow : out std_logic;  en_adder : in std_logic);
   end component;
   
   component logic_op_unit_Nbit32
      port( op1, op2 : in std_logic_vector (31 downto 0);  en_logic, s3, s2, s1
            , s0 : in std_logic;  logic_out : out std_logic_vector (31 downto 
            0));
   end component;
   
   component ALU_decoder
      port( s5, s4, s3, s2, s1, s0, en_ALU : in std_logic;  en_mult, en_comp, 
            en_Shift, en_Adder, en_Logic : out std_logic);
   end component;
   
   signal en_mult, en_comp, en_Shift, en_Adder, en_logic, out_logic_31_port, 
      out_logic_30_port, out_logic_29_port, out_logic_28_port, 
      out_logic_27_port, out_logic_26_port, out_logic_25_port, 
      out_logic_24_port, out_logic_23_port, out_logic_22_port, 
      out_logic_21_port, out_logic_20_port, out_logic_19_port, 
      out_logic_18_port, out_logic_17_port, out_logic_16_port, 
      out_logic_15_port, out_logic_14_port, out_logic_13_port, 
      out_logic_12_port, out_logic_11_port, out_logic_10_port, out_logic_9_port
      , out_logic_8_port, out_logic_7_port, out_logic_6_port, out_logic_5_port,
      out_logic_4_port, out_logic_3_port, out_logic_2_port, out_logic_1_port, 
      out_logic_0_port, out_add_31_port, out_add_30_port, out_add_29_port, 
      out_add_28_port, out_add_27_port, out_add_26_port, out_add_25_port, 
      out_add_24_port, out_add_23_port, out_add_22_port, out_add_21_port, 
      out_add_20_port, out_add_19_port, out_add_18_port, out_add_17_port, 
      out_add_16_port, out_add_15_port, out_add_14_port, out_add_13_port, 
      out_add_12_port, out_add_11_port, out_add_10_port, out_add_9_port, 
      out_add_8_port, out_add_7_port, out_add_6_port, out_add_5_port, 
      out_add_4_port, out_add_3_port, out_add_2_port, out_add_1_port, 
      out_add_0_port, out_mul_31_port, out_mul_30_port, out_mul_29_port, 
      out_mul_28_port, out_mul_27_port, out_mul_26_port, out_mul_25_port, 
      out_mul_24_port, out_mul_23_port, out_mul_22_port, out_mul_21_port, 
      out_mul_20_port, out_mul_19_port, out_mul_18_port, out_mul_17_port, 
      out_mul_16_port, out_mul_15_port, out_mul_14_port, out_mul_13_port, 
      out_mul_12_port, out_mul_11_port, out_mul_10_port, out_mul_9_port, 
      out_mul_8_port, out_mul_7_port, out_mul_6_port, out_mul_5_port, 
      out_mul_4_port, out_mul_3_port, out_mul_2_port, out_mul_1_port, 
      out_mul_0_port, out_comp_9_port, out_shift_31_port, out_shift_30_port, 
      out_shift_29_port, out_shift_28_port, out_shift_27_port, 
      out_shift_26_port, out_shift_25_port, out_shift_24_port, 
      out_shift_23_port, out_shift_22_port, out_shift_21_port, 
      out_shift_20_port, out_shift_19_port, out_shift_18_port, 
      out_shift_17_port, out_shift_16_port, out_shift_15_port, 
      out_shift_14_port, out_shift_13_port, out_shift_12_port, 
      out_shift_11_port, out_shift_10_port, out_shift_9_port, out_shift_8_port,
      out_shift_7_port, out_shift_6_port, out_shift_5_port, out_shift_4_port, 
      out_shift_3_port, out_shift_2_port, out_shift_1_port, out_shift_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n_1431
      , n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440,
      n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, 
      n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, 
      n_1459, n_1460, n_1461, n_1462, n_1463 : std_logic;

begin
   
   decoder : ALU_decoder port map( s5 => sel(5), s4 => sel(4), s3 => sel(3), s2
                           => sel(2), s1 => sel(1), s0 => sel(0), en_ALU => 
                           en_alu, en_mult => en_mult, en_comp => en_comp, 
                           en_Shift => en_Shift, en_Adder => en_Adder, en_Logic
                           => en_logic);
   logic_op : logic_op_unit_Nbit32 port map( op1(31) => op1(31), op1(30) => 
                           op1(30), op1(29) => op1(29), op1(28) => op1(28), 
                           op1(27) => op1(27), op1(26) => op1(26), op1(25) => 
                           op1(25), op1(24) => op1(24), op1(23) => op1(23), 
                           op1(22) => op1(22), op1(21) => op1(21), op1(20) => 
                           op1(20), op1(19) => op1(19), op1(18) => op1(18), 
                           op1(17) => op1(17), op1(16) => op1(16), op1(15) => 
                           n1, op1(14) => op1(14), op1(13) => op1(13), op1(12) 
                           => op1(12), op1(11) => op1(11), op1(10) => op1(10), 
                           op1(9) => op1(9), op1(8) => op1(8), op1(7) => op1(7)
                           , op1(6) => op1(6), op1(5) => op1(5), op1(4) => 
                           op1(4), op1(3) => op1(3), op1(2) => op1(2), op1(1) 
                           => op1(1), op1(0) => op1(0), op2(31) => op2(31), 
                           op2(30) => op2(30), op2(29) => op2(29), op2(28) => 
                           op2(28), op2(27) => op2(27), op2(26) => op2(26), 
                           op2(25) => op2(25), op2(24) => op2(24), op2(23) => 
                           op2(23), op2(22) => op2(22), op2(21) => op2(21), 
                           op2(20) => op2(20), op2(19) => op2(19), op2(18) => 
                           op2(18), op2(17) => op2(17), op2(16) => op2(16), 
                           op2(15) => op2(15), op2(14) => op2(14), op2(13) => 
                           op2(13), op2(12) => op2(12), op2(11) => op2(11), 
                           op2(10) => op2(10), op2(9) => op2(9), op2(8) => 
                           op2(8), op2(7) => op2(7), op2(6) => op2(6), op2(5) 
                           => op2(5), op2(4) => op2(4), op2(3) => op2(3), 
                           op2(2) => op2(2), op2(1) => op2(1), op2(0) => op2(0)
                           , en_logic => en_logic, s3 => sel(3), s2 => sel(2), 
                           s1 => sel(1), s0 => sel(0), logic_out(31) => 
                           out_logic_31_port, logic_out(30) => 
                           out_logic_30_port, logic_out(29) => 
                           out_logic_29_port, logic_out(28) => 
                           out_logic_28_port, logic_out(27) => 
                           out_logic_27_port, logic_out(26) => 
                           out_logic_26_port, logic_out(25) => 
                           out_logic_25_port, logic_out(24) => 
                           out_logic_24_port, logic_out(23) => 
                           out_logic_23_port, logic_out(22) => 
                           out_logic_22_port, logic_out(21) => 
                           out_logic_21_port, logic_out(20) => 
                           out_logic_20_port, logic_out(19) => 
                           out_logic_19_port, logic_out(18) => 
                           out_logic_18_port, logic_out(17) => 
                           out_logic_17_port, logic_out(16) => 
                           out_logic_16_port, logic_out(15) => 
                           out_logic_15_port, logic_out(14) => 
                           out_logic_14_port, logic_out(13) => 
                           out_logic_13_port, logic_out(12) => 
                           out_logic_12_port, logic_out(11) => 
                           out_logic_11_port, logic_out(10) => 
                           out_logic_10_port, logic_out(9) => out_logic_9_port,
                           logic_out(8) => out_logic_8_port, logic_out(7) => 
                           out_logic_7_port, logic_out(6) => out_logic_6_port, 
                           logic_out(5) => out_logic_5_port, logic_out(4) => 
                           out_logic_4_port, logic_out(3) => out_logic_3_port, 
                           logic_out(2) => out_logic_2_port, logic_out(1) => 
                           out_logic_1_port, logic_out(0) => out_logic_0_port);
   add_sub : adder_wrapper_nbit32 port map( op1(31) => op1(31), op1(30) => 
                           op1(30), op1(29) => op1(29), op1(28) => op1(28), 
                           op1(27) => op1(27), op1(26) => op1(26), op1(25) => 
                           op1(25), op1(24) => op1(24), op1(23) => op1(23), 
                           op1(22) => op1(22), op1(21) => op1(21), op1(20) => 
                           op1(20), op1(19) => op1(19), op1(18) => op1(18), 
                           op1(17) => op1(17), op1(16) => op1(16), op1(15) => 
                           n1, op1(14) => op1(14), op1(13) => op1(13), op1(12) 
                           => op1(12), op1(11) => op1(11), op1(10) => op1(10), 
                           op1(9) => op1(9), op1(8) => op1(8), op1(7) => op1(7)
                           , op1(6) => op1(6), op1(5) => op1(5), op1(4) => 
                           op1(4), op1(3) => op1(3), op1(2) => op1(2), op1(1) 
                           => op1(1), op1(0) => op1(0), op2(31) => op2(31), 
                           op2(30) => op2(30), op2(29) => op2(29), op2(28) => 
                           op2(28), op2(27) => op2(27), op2(26) => op2(26), 
                           op2(25) => op2(25), op2(24) => op2(24), op2(23) => 
                           op2(23), op2(22) => op2(22), op2(21) => op2(21), 
                           op2(20) => op2(20), op2(19) => op2(19), op2(18) => 
                           op2(18), op2(17) => op2(17), op2(16) => op2(16), 
                           op2(15) => op2(15), op2(14) => op2(14), op2(13) => 
                           op2(13), op2(12) => op2(12), op2(11) => op2(11), 
                           op2(10) => op2(10), op2(9) => op2(9), op2(8) => 
                           op2(8), op2(7) => op2(7), op2(6) => op2(6), op2(5) 
                           => op2(5), op2(4) => op2(4), op2(3) => op2(3), 
                           op2(2) => op2(2), op2(1) => op2(1), op2(0) => op2(0)
                           , CarryIn => sel(0), sum(31) => out_add_31_port, 
                           sum(30) => out_add_30_port, sum(29) => 
                           out_add_29_port, sum(28) => out_add_28_port, sum(27)
                           => out_add_27_port, sum(26) => out_add_26_port, 
                           sum(25) => out_add_25_port, sum(24) => 
                           out_add_24_port, sum(23) => out_add_23_port, sum(22)
                           => out_add_22_port, sum(21) => out_add_21_port, 
                           sum(20) => out_add_20_port, sum(19) => 
                           out_add_19_port, sum(18) => out_add_18_port, sum(17)
                           => out_add_17_port, sum(16) => out_add_16_port, 
                           sum(15) => out_add_15_port, sum(14) => 
                           out_add_14_port, sum(13) => out_add_13_port, sum(12)
                           => out_add_12_port, sum(11) => out_add_11_port, 
                           sum(10) => out_add_10_port, sum(9) => out_add_9_port
                           , sum(8) => out_add_8_port, sum(7) => out_add_7_port
                           , sum(6) => out_add_6_port, sum(5) => out_add_5_port
                           , sum(4) => out_add_4_port, sum(3) => out_add_3_port
                           , sum(2) => out_add_2_port, sum(1) => out_add_1_port
                           , sum(0) => out_add_0_port, CarryOut => n_1431, 
                           overflow => n_1432, en_adder => en_Adder);
   mul : mul_wrapper_NBIT32_N16_M16 port map( a(31) => op1(31), a(30) => 
                           op1(30), a(29) => op1(29), a(28) => op1(28), a(27) 
                           => op1(27), a(26) => op1(26), a(25) => op1(25), 
                           a(24) => op1(24), a(23) => op1(23), a(22) => op1(22)
                           , a(21) => op1(21), a(20) => op1(20), a(19) => 
                           op1(19), a(18) => op1(18), a(17) => op1(17), a(16) 
                           => op1(16), a(15) => n1, a(14) => op1(14), a(13) => 
                           op1(13), a(12) => op1(12), a(11) => op1(11), a(10) 
                           => op1(10), a(9) => op1(9), a(8) => op1(8), a(7) => 
                           op1(7), a(6) => op1(6), a(5) => op1(5), a(4) => 
                           op1(4), a(3) => op1(3), a(2) => op1(2), a(1) => 
                           op1(1), a(0) => op1(0), b(31) => op2(31), b(30) => 
                           op2(30), b(29) => op2(29), b(28) => op2(28), b(27) 
                           => op2(27), b(26) => op2(26), b(25) => op2(25), 
                           b(24) => op2(24), b(23) => op2(23), b(22) => op2(22)
                           , b(21) => op2(21), b(20) => op2(20), b(19) => 
                           op2(19), b(18) => op2(18), b(17) => op2(17), b(16) 
                           => op2(16), b(15) => op2(15), b(14) => op2(14), 
                           b(13) => op2(13), b(12) => op2(12), b(11) => op2(11)
                           , b(10) => op2(10), b(9) => op2(9), b(8) => op2(8), 
                           b(7) => op2(7), b(6) => op2(6), b(5) => op2(5), b(4)
                           => op2(4), b(3) => op2(3), b(2) => op2(2), b(1) => 
                           op2(1), b(0) => op2(0), en => en_mult, mul(31) => 
                           out_mul_31_port, mul(30) => out_mul_30_port, mul(29)
                           => out_mul_29_port, mul(28) => out_mul_28_port, 
                           mul(27) => out_mul_27_port, mul(26) => 
                           out_mul_26_port, mul(25) => out_mul_25_port, mul(24)
                           => out_mul_24_port, mul(23) => out_mul_23_port, 
                           mul(22) => out_mul_22_port, mul(21) => 
                           out_mul_21_port, mul(20) => out_mul_20_port, mul(19)
                           => out_mul_19_port, mul(18) => out_mul_18_port, 
                           mul(17) => out_mul_17_port, mul(16) => 
                           out_mul_16_port, mul(15) => out_mul_15_port, mul(14)
                           => out_mul_14_port, mul(13) => out_mul_13_port, 
                           mul(12) => out_mul_12_port, mul(11) => 
                           out_mul_11_port, mul(10) => out_mul_10_port, mul(9) 
                           => out_mul_9_port, mul(8) => out_mul_8_port, mul(7) 
                           => out_mul_7_port, mul(6) => out_mul_6_port, mul(5) 
                           => out_mul_5_port, mul(4) => out_mul_4_port, mul(3) 
                           => out_mul_3_port, mul(2) => out_mul_2_port, mul(1) 
                           => out_mul_1_port, mul(0) => out_mul_0_port);
   comp : zero_comparator_N32 port map( A(31) => op1(31), A(30) => op1(30), 
                           A(29) => op1(29), A(28) => op1(28), A(27) => op1(27)
                           , A(26) => op1(26), A(25) => op1(25), A(24) => 
                           op1(24), A(23) => op1(23), A(22) => op1(22), A(21) 
                           => op1(21), A(20) => op1(20), A(19) => op1(19), 
                           A(18) => op1(18), A(17) => op1(17), A(16) => op1(16)
                           , A(15) => n1, A(14) => op1(14), A(13) => op1(13), 
                           A(12) => op1(12), A(11) => op1(11), A(10) => op1(10)
                           , A(9) => op1(9), A(8) => op1(8), A(7) => op1(7), 
                           A(6) => op1(6), A(5) => op1(5), A(4) => op1(4), A(3)
                           => op1(3), A(2) => op1(2), A(1) => op1(1), A(0) => 
                           op1(0), B(31) => op2(31), B(30) => op2(30), B(29) =>
                           op2(29), B(28) => op2(28), B(27) => op2(27), B(26) 
                           => op2(26), B(25) => op2(25), B(24) => op2(24), 
                           B(23) => op2(23), B(22) => op2(22), B(21) => op2(21)
                           , B(20) => op2(20), B(19) => op2(19), B(18) => 
                           op2(18), B(17) => op2(17), B(16) => op2(16), B(15) 
                           => op2(15), B(14) => op2(14), B(13) => op2(13), 
                           B(12) => op2(12), B(11) => op2(11), B(10) => op2(10)
                           , B(9) => op2(9), B(8) => op2(8), B(7) => op2(7), 
                           B(6) => op2(6), B(5) => op2(5), B(4) => op2(4), B(3)
                           => op2(3), B(2) => op2(2), B(1) => op2(1), B(0) => 
                           op2(0), en => en_comp, cond(2) => sel(2), cond(1) =>
                           sel(1), cond(0) => sel(0), O(31) => n_1433, O(30) =>
                           n_1434, O(29) => n_1435, O(28) => n_1436, O(27) => 
                           n_1437, O(26) => n_1438, O(25) => n_1439, O(24) => 
                           n_1440, O(23) => n_1441, O(22) => n_1442, O(21) => 
                           n_1443, O(20) => n_1444, O(19) => n_1445, O(18) => 
                           n_1446, O(17) => n_1447, O(16) => n_1448, O(15) => 
                           n_1449, O(14) => n_1450, O(13) => n_1451, O(12) => 
                           n_1452, O(11) => n_1453, O(10) => n_1454, O(9) => 
                           out_comp_9_port, O(8) => n_1455, O(7) => n_1456, 
                           O(6) => n_1457, O(5) => n_1458, O(4) => n_1459, O(3)
                           => n_1460, O(2) => n_1461, O(1) => n_1462, O(0) => 
                           n_1463);
   shift : shifter_wrapper_nbit32 port map( r1(31) => op1(31), r1(30) => 
                           op1(30), r1(29) => op1(29), r1(28) => op1(28), 
                           r1(27) => op1(27), r1(26) => op1(26), r1(25) => 
                           op1(25), r1(24) => op1(24), r1(23) => op1(23), 
                           r1(22) => op1(22), r1(21) => op1(21), r1(20) => 
                           op1(20), r1(19) => op1(19), r1(18) => op1(18), 
                           r1(17) => op1(17), r1(16) => op1(16), r1(15) => n1, 
                           r1(14) => op1(14), r1(13) => op1(13), r1(12) => 
                           op1(12), r1(11) => op1(11), r1(10) => op1(10), r1(9)
                           => op1(9), r1(8) => op1(8), r1(7) => op1(7), r1(6) 
                           => op1(6), r1(5) => op1(5), r1(4) => op1(4), r1(3) 
                           => op1(3), r1(2) => op1(2), r1(1) => op1(1), r1(0) 
                           => op1(0), r2(31) => op2(31), r2(30) => op2(30), 
                           r2(29) => op2(29), r2(28) => op2(28), r2(27) => 
                           op2(27), r2(26) => op2(26), r2(25) => op2(25), 
                           r2(24) => op2(24), r2(23) => op2(23), r2(22) => 
                           op2(22), r2(21) => op2(21), r2(20) => op2(20), 
                           r2(19) => op2(19), r2(18) => op2(18), r2(17) => 
                           op2(17), r2(16) => op2(16), r2(15) => op2(15), 
                           r2(14) => op2(14), r2(13) => op2(13), r2(12) => 
                           op2(12), r2(11) => op2(11), r2(10) => op2(10), r2(9)
                           => op2(9), r2(8) => op2(8), r2(7) => op2(7), r2(6) 
                           => op2(6), r2(5) => op2(5), r2(4) => op2(4), r2(3) 
                           => op2(3), r2(2) => op2(2), r2(1) => op2(1), r2(0) 
                           => op2(0), conf(1) => sel(1), conf(0) => sel(0), 
                           en_shifter => en_Shift, shifted_out(31) => 
                           out_shift_31_port, shifted_out(30) => 
                           out_shift_30_port, shifted_out(29) => 
                           out_shift_29_port, shifted_out(28) => 
                           out_shift_28_port, shifted_out(27) => 
                           out_shift_27_port, shifted_out(26) => 
                           out_shift_26_port, shifted_out(25) => 
                           out_shift_25_port, shifted_out(24) => 
                           out_shift_24_port, shifted_out(23) => 
                           out_shift_23_port, shifted_out(22) => 
                           out_shift_22_port, shifted_out(21) => 
                           out_shift_21_port, shifted_out(20) => 
                           out_shift_20_port, shifted_out(19) => 
                           out_shift_19_port, shifted_out(18) => 
                           out_shift_18_port, shifted_out(17) => 
                           out_shift_17_port, shifted_out(16) => 
                           out_shift_16_port, shifted_out(15) => 
                           out_shift_15_port, shifted_out(14) => 
                           out_shift_14_port, shifted_out(13) => 
                           out_shift_13_port, shifted_out(12) => 
                           out_shift_12_port, shifted_out(11) => 
                           out_shift_11_port, shifted_out(10) => 
                           out_shift_10_port, shifted_out(9) => 
                           out_shift_9_port, shifted_out(8) => out_shift_8_port
                           , shifted_out(7) => out_shift_7_port, shifted_out(6)
                           => out_shift_6_port, shifted_out(5) => 
                           out_shift_5_port, shifted_out(4) => out_shift_4_port
                           , shifted_out(3) => out_shift_3_port, shifted_out(2)
                           => out_shift_2_port, shifted_out(1) => 
                           out_shift_1_port, shifted_out(0) => out_shift_0_port
                           );
   U2 : AND3_X2 port map( A1 => en_comp, A2 => n70, A3 => out_comp_9_port, ZN 
                           => n6);
   U3 : AND4_X2 port map( A1 => en_logic, A2 => n71, A3 => n73, A4 => n72, ZN 
                           => n4);
   U4 : AND2_X2 port map( A1 => en_Shift, A2 => n71, ZN => n7);
   U5 : AND3_X2 port map( A1 => n71, A2 => n72, A3 => en_Adder, ZN => n5);
   U6 : BUF_X2 port map( A => op1(15), Z => n1);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => result(9));
   U8 : AOI221_X1 port map( B1 => out_logic_9_port, B2 => n4, C1 => 
                           out_add_9_port, C2 => n5, A => n6, ZN => n3);
   U9 : AOI22_X1 port map( A1 => out_shift_9_port, A2 => n7, B1 => 
                           out_mul_9_port, B2 => en_mult, ZN => n2);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => result(8));
   U11 : AOI221_X1 port map( B1 => out_logic_8_port, B2 => n4, C1 => 
                           out_add_8_port, C2 => n5, A => n6, ZN => n9);
   U12 : AOI22_X1 port map( A1 => out_shift_8_port, A2 => n7, B1 => 
                           out_mul_8_port, B2 => en_mult, ZN => n8);
   U13 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => result(7));
   U14 : AOI221_X1 port map( B1 => out_logic_7_port, B2 => n4, C1 => 
                           out_add_7_port, C2 => n5, A => n6, ZN => n11);
   U15 : AOI22_X1 port map( A1 => out_shift_7_port, A2 => n7, B1 => 
                           out_mul_7_port, B2 => en_mult, ZN => n10);
   U16 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => result(6));
   U17 : AOI221_X1 port map( B1 => out_logic_6_port, B2 => n4, C1 => 
                           out_add_6_port, C2 => n5, A => n6, ZN => n13);
   U18 : AOI22_X1 port map( A1 => out_shift_6_port, A2 => n7, B1 => 
                           out_mul_6_port, B2 => en_mult, ZN => n12);
   U19 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => result(5));
   U20 : AOI221_X1 port map( B1 => out_logic_5_port, B2 => n4, C1 => 
                           out_add_5_port, C2 => n5, A => n6, ZN => n15);
   U21 : AOI22_X1 port map( A1 => out_shift_5_port, A2 => n7, B1 => 
                           out_mul_5_port, B2 => en_mult, ZN => n14);
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => result(4));
   U23 : AOI221_X1 port map( B1 => out_logic_4_port, B2 => n4, C1 => 
                           out_add_4_port, C2 => n5, A => n6, ZN => n17);
   U24 : AOI22_X1 port map( A1 => out_shift_4_port, A2 => n7, B1 => 
                           out_mul_4_port, B2 => en_mult, ZN => n16);
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => result(3));
   U26 : AOI221_X1 port map( B1 => out_logic_3_port, B2 => n4, C1 => 
                           out_add_3_port, C2 => n5, A => n6, ZN => n19);
   U27 : AOI22_X1 port map( A1 => out_shift_3_port, A2 => n7, B1 => 
                           out_mul_3_port, B2 => en_mult, ZN => n18);
   U28 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => result(31));
   U29 : AOI221_X1 port map( B1 => out_logic_31_port, B2 => n4, C1 => 
                           out_add_31_port, C2 => n5, A => n6, ZN => n21);
   U30 : AOI22_X1 port map( A1 => out_shift_31_port, A2 => n7, B1 => 
                           out_mul_31_port, B2 => en_mult, ZN => n20);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => result(30));
   U32 : AOI221_X1 port map( B1 => out_logic_30_port, B2 => n4, C1 => 
                           out_add_30_port, C2 => n5, A => n6, ZN => n23);
   U33 : AOI22_X1 port map( A1 => out_shift_30_port, A2 => n7, B1 => 
                           out_mul_30_port, B2 => en_mult, ZN => n22);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => result(2));
   U35 : AOI221_X1 port map( B1 => out_logic_2_port, B2 => n4, C1 => 
                           out_add_2_port, C2 => n5, A => n6, ZN => n25);
   U36 : AOI22_X1 port map( A1 => out_shift_2_port, A2 => n7, B1 => 
                           out_mul_2_port, B2 => en_mult, ZN => n24);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => result(29));
   U38 : AOI221_X1 port map( B1 => out_logic_29_port, B2 => n4, C1 => 
                           out_add_29_port, C2 => n5, A => n6, ZN => n27);
   U39 : AOI22_X1 port map( A1 => out_shift_29_port, A2 => n7, B1 => 
                           out_mul_29_port, B2 => en_mult, ZN => n26);
   U40 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => result(28));
   U41 : AOI221_X1 port map( B1 => out_logic_28_port, B2 => n4, C1 => 
                           out_add_28_port, C2 => n5, A => n6, ZN => n29);
   U42 : AOI22_X1 port map( A1 => out_shift_28_port, A2 => n7, B1 => 
                           out_mul_28_port, B2 => en_mult, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => result(27));
   U44 : AOI221_X1 port map( B1 => out_logic_27_port, B2 => n4, C1 => 
                           out_add_27_port, C2 => n5, A => n6, ZN => n31);
   U45 : AOI22_X1 port map( A1 => out_shift_27_port, A2 => n7, B1 => 
                           out_mul_27_port, B2 => en_mult, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => result(26));
   U47 : AOI221_X1 port map( B1 => out_logic_26_port, B2 => n4, C1 => 
                           out_add_26_port, C2 => n5, A => n6, ZN => n33);
   U48 : AOI22_X1 port map( A1 => out_shift_26_port, A2 => n7, B1 => 
                           out_mul_26_port, B2 => en_mult, ZN => n32);
   U49 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => result(25));
   U50 : AOI221_X1 port map( B1 => out_logic_25_port, B2 => n4, C1 => 
                           out_add_25_port, C2 => n5, A => n6, ZN => n35);
   U51 : AOI22_X1 port map( A1 => out_shift_25_port, A2 => n7, B1 => 
                           out_mul_25_port, B2 => en_mult, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => result(24));
   U53 : AOI221_X1 port map( B1 => out_logic_24_port, B2 => n4, C1 => 
                           out_add_24_port, C2 => n5, A => n6, ZN => n37);
   U54 : AOI22_X1 port map( A1 => out_shift_24_port, A2 => n7, B1 => 
                           out_mul_24_port, B2 => en_mult, ZN => n36);
   U55 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => result(23));
   U56 : AOI221_X1 port map( B1 => out_logic_23_port, B2 => n4, C1 => 
                           out_add_23_port, C2 => n5, A => n6, ZN => n39);
   U57 : AOI22_X1 port map( A1 => out_shift_23_port, A2 => n7, B1 => 
                           out_mul_23_port, B2 => en_mult, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => result(22));
   U59 : AOI221_X1 port map( B1 => out_logic_22_port, B2 => n4, C1 => 
                           out_add_22_port, C2 => n5, A => n6, ZN => n41);
   U60 : AOI22_X1 port map( A1 => out_shift_22_port, A2 => n7, B1 => 
                           out_mul_22_port, B2 => en_mult, ZN => n40);
   U61 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => result(21));
   U62 : AOI221_X1 port map( B1 => out_logic_21_port, B2 => n4, C1 => 
                           out_add_21_port, C2 => n5, A => n6, ZN => n43);
   U63 : AOI22_X1 port map( A1 => out_shift_21_port, A2 => n7, B1 => 
                           out_mul_21_port, B2 => en_mult, ZN => n42);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => result(20));
   U65 : AOI221_X1 port map( B1 => out_logic_20_port, B2 => n4, C1 => 
                           out_add_20_port, C2 => n5, A => n6, ZN => n45);
   U66 : AOI22_X1 port map( A1 => out_shift_20_port, A2 => n7, B1 => 
                           out_mul_20_port, B2 => en_mult, ZN => n44);
   U67 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => result(1));
   U68 : AOI221_X1 port map( B1 => out_logic_1_port, B2 => n4, C1 => 
                           out_add_1_port, C2 => n5, A => n6, ZN => n47);
   U69 : AOI22_X1 port map( A1 => out_shift_1_port, A2 => n7, B1 => 
                           out_mul_1_port, B2 => en_mult, ZN => n46);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => result(19));
   U71 : AOI221_X1 port map( B1 => out_logic_19_port, B2 => n4, C1 => 
                           out_add_19_port, C2 => n5, A => n6, ZN => n49);
   U72 : AOI22_X1 port map( A1 => out_shift_19_port, A2 => n7, B1 => 
                           out_mul_19_port, B2 => en_mult, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => result(18));
   U74 : AOI221_X1 port map( B1 => out_logic_18_port, B2 => n4, C1 => 
                           out_add_18_port, C2 => n5, A => n6, ZN => n51);
   U75 : AOI22_X1 port map( A1 => out_shift_18_port, A2 => n7, B1 => 
                           out_mul_18_port, B2 => en_mult, ZN => n50);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => result(17));
   U77 : AOI221_X1 port map( B1 => out_logic_17_port, B2 => n4, C1 => 
                           out_add_17_port, C2 => n5, A => n6, ZN => n53);
   U78 : AOI22_X1 port map( A1 => out_shift_17_port, A2 => n7, B1 => 
                           out_mul_17_port, B2 => en_mult, ZN => n52);
   U79 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => result(16));
   U80 : AOI221_X1 port map( B1 => out_logic_16_port, B2 => n4, C1 => 
                           out_add_16_port, C2 => n5, A => n6, ZN => n55);
   U81 : AOI22_X1 port map( A1 => out_shift_16_port, A2 => n7, B1 => 
                           out_mul_16_port, B2 => en_mult, ZN => n54);
   U82 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => result(15));
   U83 : AOI221_X1 port map( B1 => out_logic_15_port, B2 => n4, C1 => 
                           out_add_15_port, C2 => n5, A => n6, ZN => n57);
   U84 : AOI22_X1 port map( A1 => out_shift_15_port, A2 => n7, B1 => 
                           out_mul_15_port, B2 => en_mult, ZN => n56);
   U85 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => result(14));
   U86 : AOI221_X1 port map( B1 => out_logic_14_port, B2 => n4, C1 => 
                           out_add_14_port, C2 => n5, A => n6, ZN => n59);
   U87 : AOI22_X1 port map( A1 => out_shift_14_port, A2 => n7, B1 => 
                           out_mul_14_port, B2 => en_mult, ZN => n58);
   U88 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => result(13));
   U89 : AOI221_X1 port map( B1 => out_logic_13_port, B2 => n4, C1 => 
                           out_add_13_port, C2 => n5, A => n6, ZN => n61);
   U90 : AOI22_X1 port map( A1 => out_shift_13_port, A2 => n7, B1 => 
                           out_mul_13_port, B2 => en_mult, ZN => n60);
   U91 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => result(12));
   U92 : AOI221_X1 port map( B1 => out_logic_12_port, B2 => n4, C1 => 
                           out_add_12_port, C2 => n5, A => n6, ZN => n63);
   U93 : AOI22_X1 port map( A1 => out_shift_12_port, A2 => n7, B1 => 
                           out_mul_12_port, B2 => en_mult, ZN => n62);
   U94 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => result(11));
   U95 : AOI221_X1 port map( B1 => out_logic_11_port, B2 => n4, C1 => 
                           out_add_11_port, C2 => n5, A => n6, ZN => n65);
   U96 : AOI22_X1 port map( A1 => out_shift_11_port, A2 => n7, B1 => 
                           out_mul_11_port, B2 => en_mult, ZN => n64);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => result(10));
   U98 : AOI221_X1 port map( B1 => out_logic_10_port, B2 => n4, C1 => 
                           out_add_10_port, C2 => n5, A => n6, ZN => n67);
   U99 : AOI22_X1 port map( A1 => out_shift_10_port, A2 => n7, B1 => 
                           out_mul_10_port, B2 => en_mult, ZN => n66);
   U100 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => result(0));
   U101 : AOI221_X1 port map( B1 => out_logic_0_port, B2 => n4, C1 => 
                           out_add_0_port, C2 => n5, A => n6, ZN => n69);
   U102 : INV_X1 port map( A => en_mult, ZN => n70);
   U103 : INV_X1 port map( A => en_Shift, ZN => n72);
   U104 : INV_X1 port map( A => en_Adder, ZN => n73);
   U105 : AOI22_X1 port map( A1 => out_shift_0_port, A2 => n7, B1 => 
                           out_mul_0_port, B2 => en_mult, ZN => n68);
   U106 : NOR2_X1 port map( A1 => en_comp, A2 => en_mult, ZN => n71);

end SYN_Specification;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity mux31_N32_0 is

   port( a, b, c : in std_logic_vector (31 downto 0);  sel : in 
         std_logic_vector (1 downto 0);  y : out std_logic_vector (31 downto 0)
         );

end mux31_N32_0;

architecture SYN_Behavioral of mux31_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X2
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n72, N37, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37_port, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : 
      std_logic;

begin
   
   y_reg_31_inst : DLH_X1 port map( G => N37, D => n71, Q => y(31));
   y_reg_30_inst : DLH_X1 port map( G => N37, D => n70, Q => y(30));
   y_reg_29_inst : DLH_X1 port map( G => N37, D => n69, Q => y(29));
   y_reg_28_inst : DLH_X1 port map( G => N37, D => n68, Q => y(28));
   y_reg_27_inst : DLH_X1 port map( G => N37, D => n67, Q => y(27));
   y_reg_26_inst : DLH_X1 port map( G => N37, D => n66, Q => y(26));
   y_reg_25_inst : DLH_X1 port map( G => N37, D => n65, Q => y(25));
   y_reg_24_inst : DLH_X1 port map( G => N37, D => n64, Q => y(24));
   y_reg_23_inst : DLH_X1 port map( G => N37, D => n63, Q => y(23));
   y_reg_22_inst : DLH_X1 port map( G => N37, D => n62, Q => y(22));
   y_reg_21_inst : DLH_X1 port map( G => N37, D => n61, Q => y(21));
   y_reg_20_inst : DLH_X1 port map( G => N37, D => n60, Q => y(20));
   y_reg_19_inst : DLH_X1 port map( G => N37, D => n59, Q => y(19));
   y_reg_18_inst : DLH_X1 port map( G => N37, D => n58, Q => y(18));
   y_reg_17_inst : DLH_X1 port map( G => N37, D => n57, Q => y(17));
   y_reg_16_inst : DLH_X1 port map( G => N37, D => n56, Q => y(16));
   y_reg_15_inst : DLH_X1 port map( G => N37, D => n55, Q => y(15));
   y_reg_0_inst : DLH_X1 port map( G => N37, D => n40, Q => n72);
   y_reg_1_inst : DLH_X2 port map( G => N37, D => n41, Q => y(1));
   y_reg_9_inst : DLH_X2 port map( G => N37, D => n49, Q => y(9));
   y_reg_12_inst : DLH_X2 port map( G => N37, D => n52, Q => y(12));
   y_reg_5_inst : DLH_X2 port map( G => N37, D => n45, Q => y(5));
   y_reg_8_inst : DLH_X2 port map( G => N37, D => n48, Q => y(8));
   y_reg_11_inst : DLH_X2 port map( G => N37, D => n51, Q => y(11));
   y_reg_4_inst : DLH_X2 port map( G => N37, D => n44, Q => y(4));
   y_reg_2_inst : DLH_X2 port map( G => N37, D => n42, Q => y(2));
   y_reg_14_inst : DLH_X2 port map( G => N37, D => n54, Q => y(14));
   y_reg_10_inst : DLH_X2 port map( G => N37, D => n50, Q => y(10));
   y_reg_7_inst : DLH_X2 port map( G => N37, D => n47, Q => y(7));
   y_reg_3_inst : DLH_X2 port map( G => N37, D => n43, Q => y(3));
   y_reg_13_inst : DLH_X2 port map( G => N37, D => n53, Q => y(13));
   y_reg_6_inst : DLH_X2 port map( G => N37, D => n46, Q => y(6));
   U3 : OR2_X1 port map( A1 => n3, A2 => n7, ZN => n1);
   U4 : OR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n2);
   U5 : INV_X2 port map( A => n2, ZN => n3);
   U6 : INV_X2 port map( A => n1, ZN => n4);
   U7 : CLKBUF_X3 port map( A => n72, Z => y(0));
   U8 : NOR2_X4 port map( A1 => n39, A2 => sel(1), ZN => n7);
   U9 : INV_X1 port map( A => n6, ZN => n40);
   U10 : AOI222_X1 port map( A1 => b(0), A2 => n7, B1 => c(0), B2 => n4, C1 => 
                           a(0), C2 => n3, ZN => n6);
   U11 : INV_X1 port map( A => n8, ZN => n41);
   U12 : AOI222_X1 port map( A1 => b(1), A2 => n7, B1 => c(1), B2 => n4, C1 => 
                           a(1), C2 => n3, ZN => n8);
   U13 : INV_X1 port map( A => n9, ZN => n42);
   U14 : AOI222_X1 port map( A1 => b(2), A2 => n7, B1 => c(2), B2 => n4, C1 => 
                           a(2), C2 => n3, ZN => n9);
   U15 : INV_X1 port map( A => n10, ZN => n43);
   U16 : AOI222_X1 port map( A1 => b(3), A2 => n7, B1 => c(3), B2 => n4, C1 => 
                           a(3), C2 => n3, ZN => n10);
   U17 : INV_X1 port map( A => n11, ZN => n44);
   U18 : AOI222_X1 port map( A1 => b(4), A2 => n7, B1 => c(4), B2 => n4, C1 => 
                           a(4), C2 => n3, ZN => n11);
   U19 : INV_X1 port map( A => n12, ZN => n45);
   U20 : AOI222_X1 port map( A1 => b(5), A2 => n7, B1 => c(5), B2 => n4, C1 => 
                           a(5), C2 => n3, ZN => n12);
   U21 : INV_X1 port map( A => n13, ZN => n46);
   U22 : AOI222_X1 port map( A1 => b(6), A2 => n7, B1 => c(6), B2 => n4, C1 => 
                           a(6), C2 => n3, ZN => n13);
   U23 : INV_X1 port map( A => n14, ZN => n47);
   U24 : AOI222_X1 port map( A1 => b(7), A2 => n7, B1 => c(7), B2 => n4, C1 => 
                           a(7), C2 => n3, ZN => n14);
   U25 : INV_X1 port map( A => n15, ZN => n48);
   U26 : AOI222_X1 port map( A1 => b(8), A2 => n7, B1 => c(8), B2 => n4, C1 => 
                           a(8), C2 => n3, ZN => n15);
   U27 : INV_X1 port map( A => n16, ZN => n49);
   U28 : AOI222_X1 port map( A1 => b(9), A2 => n7, B1 => c(9), B2 => n4, C1 => 
                           a(9), C2 => n3, ZN => n16);
   U29 : INV_X1 port map( A => n17, ZN => n50);
   U30 : AOI222_X1 port map( A1 => b(10), A2 => n7, B1 => c(10), B2 => n4, C1 
                           => a(10), C2 => n3, ZN => n17);
   U31 : INV_X1 port map( A => n18, ZN => n51);
   U32 : AOI222_X1 port map( A1 => b(11), A2 => n7, B1 => c(11), B2 => n4, C1 
                           => a(11), C2 => n3, ZN => n18);
   U33 : INV_X1 port map( A => n19, ZN => n52);
   U34 : AOI222_X1 port map( A1 => b(12), A2 => n7, B1 => c(12), B2 => n4, C1 
                           => a(12), C2 => n3, ZN => n19);
   U35 : INV_X1 port map( A => n20, ZN => n53);
   U36 : AOI222_X1 port map( A1 => b(13), A2 => n7, B1 => c(13), B2 => n4, C1 
                           => a(13), C2 => n3, ZN => n20);
   U37 : INV_X1 port map( A => n21, ZN => n54);
   U38 : AOI222_X1 port map( A1 => b(14), A2 => n7, B1 => c(14), B2 => n4, C1 
                           => a(14), C2 => n3, ZN => n21);
   U39 : INV_X1 port map( A => n22, ZN => n55);
   U40 : AOI222_X1 port map( A1 => b(15), A2 => n7, B1 => c(15), B2 => n4, C1 
                           => a(15), C2 => n3, ZN => n22);
   U41 : INV_X1 port map( A => n23, ZN => n56);
   U42 : AOI222_X1 port map( A1 => b(16), A2 => n7, B1 => c(16), B2 => n4, C1 
                           => a(16), C2 => n3, ZN => n23);
   U43 : INV_X1 port map( A => n24, ZN => n57);
   U44 : AOI222_X1 port map( A1 => b(17), A2 => n7, B1 => c(17), B2 => n4, C1 
                           => a(17), C2 => n3, ZN => n24);
   U45 : INV_X1 port map( A => n25, ZN => n58);
   U46 : AOI222_X1 port map( A1 => b(18), A2 => n7, B1 => c(18), B2 => n4, C1 
                           => a(18), C2 => n3, ZN => n25);
   U47 : INV_X1 port map( A => n26, ZN => n59);
   U48 : AOI222_X1 port map( A1 => b(19), A2 => n7, B1 => c(19), B2 => n4, C1 
                           => a(19), C2 => n3, ZN => n26);
   U49 : INV_X1 port map( A => n27, ZN => n60);
   U50 : AOI222_X1 port map( A1 => b(20), A2 => n7, B1 => c(20), B2 => n4, C1 
                           => a(20), C2 => n3, ZN => n27);
   U51 : INV_X1 port map( A => n28, ZN => n61);
   U52 : AOI222_X1 port map( A1 => b(21), A2 => n7, B1 => c(21), B2 => n4, C1 
                           => a(21), C2 => n3, ZN => n28);
   U53 : INV_X1 port map( A => n29, ZN => n62);
   U54 : AOI222_X1 port map( A1 => b(22), A2 => n7, B1 => c(22), B2 => n4, C1 
                           => a(22), C2 => n3, ZN => n29);
   U55 : INV_X1 port map( A => n30, ZN => n63);
   U56 : AOI222_X1 port map( A1 => b(23), A2 => n7, B1 => c(23), B2 => n4, C1 
                           => a(23), C2 => n3, ZN => n30);
   U57 : INV_X1 port map( A => n31, ZN => n64);
   U58 : AOI222_X1 port map( A1 => b(24), A2 => n7, B1 => c(24), B2 => n4, C1 
                           => a(24), C2 => n3, ZN => n31);
   U59 : INV_X1 port map( A => n32, ZN => n65);
   U60 : AOI222_X1 port map( A1 => b(25), A2 => n7, B1 => c(25), B2 => n4, C1 
                           => a(25), C2 => n3, ZN => n32);
   U61 : INV_X1 port map( A => n33, ZN => n66);
   U62 : AOI222_X1 port map( A1 => b(26), A2 => n7, B1 => c(26), B2 => n4, C1 
                           => a(26), C2 => n3, ZN => n33);
   U63 : INV_X1 port map( A => n34, ZN => n67);
   U64 : AOI222_X1 port map( A1 => b(27), A2 => n7, B1 => c(27), B2 => n4, C1 
                           => a(27), C2 => n3, ZN => n34);
   U65 : INV_X1 port map( A => n35, ZN => n68);
   U66 : AOI222_X1 port map( A1 => b(28), A2 => n7, B1 => c(28), B2 => n4, C1 
                           => a(28), C2 => n3, ZN => n35);
   U67 : INV_X1 port map( A => n36, ZN => n69);
   U68 : AOI222_X1 port map( A1 => b(29), A2 => n7, B1 => c(29), B2 => n4, C1 
                           => a(29), C2 => n3, ZN => n36);
   U69 : INV_X1 port map( A => n37_port, ZN => n70);
   U70 : AOI222_X1 port map( A1 => b(30), A2 => n7, B1 => c(30), B2 => n4, C1 
                           => a(30), C2 => n3, ZN => n37_port);
   U71 : INV_X1 port map( A => n38, ZN => n71);
   U72 : AOI222_X1 port map( A1 => b(31), A2 => n7, B1 => c(31), B2 => n4, C1 
                           => a(31), C2 => n3, ZN => n38);
   U73 : NAND2_X1 port map( A1 => n4, A2 => sel(0), ZN => N37);
   U74 : INV_X1 port map( A => sel(0), ZN => n39);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity comparator_addr is

   port( y1, y2 : in std_logic_vector (31 downto 0);  comp_control : in 
         std_logic_vector (1 downto 0);  EqualD : out std_logic);

end comparator_addr;

architecture SYN_Behavioral of comparator_addr is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component comparator_addr_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N6, N44, n1, n4, n2, n3, n5, n6_port, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n_1464, n_1465, n_1466, n_1467, n_1468 : std_logic;

begin
   
   n1 <= '0';
   EqualD_reg : DLH_X1 port map( G => n4, D => N44, Q => EqualD);
   n4 <= '1';
   eq_26 : comparator_addr_DW01_cmp6_0 port map( A(31) => y1(31), A(30) => 
                           y1(30), A(29) => y1(29), A(28) => y1(28), A(27) => 
                           y1(27), A(26) => y1(26), A(25) => y1(25), A(24) => 
                           y1(24), A(23) => y1(23), A(22) => y1(22), A(21) => 
                           y1(21), A(20) => y1(20), A(19) => y1(19), A(18) => 
                           y1(18), A(17) => y1(17), A(16) => y1(16), A(15) => 
                           y1(15), A(14) => y1(14), A(13) => y1(13), A(12) => 
                           y1(12), A(11) => y1(11), A(10) => y1(10), A(9) => 
                           y1(9), A(8) => y1(8), A(7) => y1(7), A(6) => y1(6), 
                           A(5) => y1(5), A(4) => y1(4), A(3) => y1(3), A(2) =>
                           y1(2), A(1) => y1(1), A(0) => y1(0), B(31) => y2(31)
                           , B(30) => y2(30), B(29) => y2(29), B(28) => y2(28),
                           B(27) => y2(27), B(26) => y2(26), B(25) => y2(25), 
                           B(24) => y2(24), B(23) => y2(23), B(22) => y2(22), 
                           B(21) => y2(21), B(20) => y2(20), B(19) => y2(19), 
                           B(18) => y2(18), B(17) => y2(17), B(16) => y2(16), 
                           B(15) => y2(15), B(14) => y2(14), B(13) => y2(13), 
                           B(12) => y2(12), B(11) => y2(11), B(10) => y2(10), 
                           B(9) => y2(9), B(8) => y2(8), B(7) => y2(7), B(6) =>
                           y2(6), B(5) => y2(5), B(4) => y2(4), B(3) => y2(3), 
                           B(2) => y2(2), B(1) => y2(1), B(0) => y2(0), TC => 
                           n1, LT => n_1464, GT => n_1465, EQ => N6, LE => 
                           n_1466, GE => n_1467, NE => n_1468);
   U3 : MUX2_X1 port map( A => n2, B => N6, S => n3, Z => N44);
   U4 : NOR2_X1 port map( A1 => comp_control(1), A2 => comp_control(0), ZN => 
                           n3);
   U6 : NAND2_X1 port map( A1 => n5, A2 => comp_control(1), ZN => n2);
   U7 : XNOR2_X1 port map( A => comp_control(0), B => n6_port, ZN => n5);
   U8 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => n6_port);
   U9 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n8)
                           ;
   U10 : NOR4_X1 port map( A1 => y1(23), A2 => y1(22), A3 => y1(21), A4 => 
                           y1(20), ZN => n12);
   U11 : NOR4_X1 port map( A1 => y1(1), A2 => y1(19), A3 => y1(18), A4 => 
                           y1(17), ZN => n11);
   U12 : NOR4_X1 port map( A1 => y1(16), A2 => y1(15), A3 => y1(14), A4 => 
                           y1(13), ZN => n10);
   U13 : NOR4_X1 port map( A1 => y1(12), A2 => y1(11), A3 => y1(10), A4 => 
                           y1(0), ZN => n9);
   U14 : NAND4_X1 port map( A1 => n13, A2 => n14, A3 => n15, A4 => n16, ZN => 
                           n7);
   U15 : NOR4_X1 port map( A1 => y1(9), A2 => y1(8), A3 => y1(7), A4 => y1(6), 
                           ZN => n16);
   U16 : NOR4_X1 port map( A1 => y1(5), A2 => y1(4), A3 => y1(3), A4 => y1(31),
                           ZN => n15);
   U17 : NOR4_X1 port map( A1 => y1(30), A2 => y1(2), A3 => y1(29), A4 => 
                           y1(28), ZN => n14);
   U18 : NOR4_X1 port map( A1 => y1(27), A2 => y1(26), A3 => y1(25), A4 => 
                           y1(24), ZN => n13);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity window_rf_M4_N4_F4_NBIT32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  WR_ADD, RD1_ADD, 
         RD2_ADD : in std_logic_vector (4 downto 0);  FILL, SPILL : out 
         std_logic;  CALL, RET : in std_logic;  MEM_IN : in std_logic_vector 
         (31 downto 0);  MEM_OUT : out std_logic_vector (31 downto 0);  DATAIN 
         : in std_logic_vector (31 downto 0);  OUT1, OUT2 : out 
         std_logic_vector (31 downto 0));

end window_rf_M4_N4_F4_NBIT32;

architecture SYN_Behavioral of window_rf_M4_N4_F4_NBIT32 is

   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X4
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component window_rf_M4_N4_F4_NBIT32_DW01_add_4
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component window_rf_M4_N4_F4_NBIT32_DW01_sub_4
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component window_rf_M4_N4_F4_NBIT32_DW01_sub_3
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component window_rf_M4_N4_F4_NBIT32_DW01_add_3
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   component window_rf_M4_N4_F4_NBIT32_DW01_add_2
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   component window_rf_M4_N4_F4_NBIT32_DW01_add_1
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   component window_rf_M4_N4_F4_NBIT32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, FILL_port, MEM_OUT_31_port, 
      MEM_OUT_30_port, MEM_OUT_29_port, MEM_OUT_28_port, MEM_OUT_27_port, 
      MEM_OUT_26_port, MEM_OUT_25_port, MEM_OUT_24_port, MEM_OUT_23_port, 
      MEM_OUT_22_port, MEM_OUT_21_port, MEM_OUT_20_port, MEM_OUT_19_port, 
      MEM_OUT_18_port, MEM_OUT_17_port, MEM_OUT_16_port, MEM_OUT_15_port, 
      MEM_OUT_14_port, MEM_OUT_13_port, MEM_OUT_12_port, MEM_OUT_11_port, 
      MEM_OUT_10_port, MEM_OUT_9_port, MEM_OUT_8_port, MEM_OUT_7_port, 
      MEM_OUT_6_port, MEM_OUT_5_port, MEM_OUT_4_port, MEM_OUT_3_port, 
      MEM_OUT_2_port, MEM_OUT_1_port, MEM_OUT_0_port, CWP_31_port, CWP_30_port,
      CWP_29_port, CWP_28_port, CWP_27_port, CWP_26_port, CWP_25_port, 
      CWP_24_port, CWP_23_port, CWP_22_port, CWP_21_port, CWP_20_port, 
      CWP_19_port, CWP_18_port, CWP_17_port, CWP_16_port, CWP_15_port, 
      CWP_14_port, CWP_13_port, CWP_12_port, CWP_11_port, CWP_10_port, 
      CWP_9_port, CWP_8_port, CWP_7_port, CWP_6_port, CWP_5_port, CWP_4_port, 
      CWP_3_port, CWP_2_port, CWP_1_port, CWP_0_port, N3564, N3565, N3566, 
      N3567, N3568, N3569, N3570, N3571, N3572, ADD_RD1_5_port, N3577, N3578, 
      N3579, N3580, N3581, N3582, N3583, N3584, N3585, ADD_RD2_5_port, N3590, 
      N3591, N3592, N3593, N3594, N3595, N3596, N3597, N3598, 
      REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, REGISTERS_32_31_port, REGISTERS_32_30_port, 
      REGISTERS_32_29_port, REGISTERS_32_28_port, REGISTERS_32_27_port, 
      REGISTERS_32_26_port, REGISTERS_32_25_port, REGISTERS_32_24_port, 
      REGISTERS_32_23_port, REGISTERS_32_22_port, REGISTERS_32_21_port, 
      REGISTERS_32_20_port, REGISTERS_32_19_port, REGISTERS_32_18_port, 
      REGISTERS_32_17_port, REGISTERS_32_16_port, REGISTERS_32_15_port, 
      REGISTERS_32_14_port, REGISTERS_32_13_port, REGISTERS_32_12_port, 
      REGISTERS_32_11_port, REGISTERS_32_10_port, REGISTERS_32_9_port, 
      REGISTERS_32_8_port, REGISTERS_32_7_port, REGISTERS_32_6_port, 
      REGISTERS_32_5_port, REGISTERS_32_4_port, REGISTERS_32_3_port, 
      REGISTERS_32_2_port, REGISTERS_32_1_port, REGISTERS_32_0_port, 
      REGISTERS_33_31_port, REGISTERS_33_30_port, REGISTERS_33_29_port, 
      REGISTERS_33_28_port, REGISTERS_33_27_port, REGISTERS_33_26_port, 
      REGISTERS_33_25_port, REGISTERS_33_24_port, REGISTERS_33_23_port, 
      REGISTERS_33_22_port, REGISTERS_33_21_port, REGISTERS_33_20_port, 
      REGISTERS_33_19_port, REGISTERS_33_18_port, REGISTERS_33_17_port, 
      REGISTERS_33_16_port, REGISTERS_33_15_port, REGISTERS_33_14_port, 
      REGISTERS_33_13_port, REGISTERS_33_12_port, REGISTERS_33_11_port, 
      REGISTERS_33_10_port, REGISTERS_33_9_port, REGISTERS_33_8_port, 
      REGISTERS_33_7_port, REGISTERS_33_6_port, REGISTERS_33_5_port, 
      REGISTERS_33_4_port, REGISTERS_33_3_port, REGISTERS_33_2_port, 
      REGISTERS_33_1_port, REGISTERS_33_0_port, REGISTERS_34_31_port, 
      REGISTERS_34_30_port, REGISTERS_34_29_port, REGISTERS_34_28_port, 
      REGISTERS_34_27_port, REGISTERS_34_26_port, REGISTERS_34_25_port, 
      REGISTERS_34_24_port, REGISTERS_34_23_port, REGISTERS_34_22_port, 
      REGISTERS_34_21_port, REGISTERS_34_20_port, REGISTERS_34_19_port, 
      REGISTERS_34_18_port, REGISTERS_34_17_port, REGISTERS_34_16_port, 
      REGISTERS_34_15_port, REGISTERS_34_14_port, REGISTERS_34_13_port, 
      REGISTERS_34_12_port, REGISTERS_34_11_port, REGISTERS_34_10_port, 
      REGISTERS_34_9_port, REGISTERS_34_8_port, REGISTERS_34_7_port, 
      REGISTERS_34_6_port, REGISTERS_34_5_port, REGISTERS_34_4_port, 
      REGISTERS_34_3_port, REGISTERS_34_2_port, REGISTERS_34_1_port, 
      REGISTERS_34_0_port, REGISTERS_35_31_port, REGISTERS_35_30_port, 
      REGISTERS_35_29_port, REGISTERS_35_28_port, REGISTERS_35_27_port, 
      REGISTERS_35_26_port, REGISTERS_35_25_port, REGISTERS_35_24_port, 
      REGISTERS_35_23_port, REGISTERS_35_22_port, REGISTERS_35_21_port, 
      REGISTERS_35_20_port, REGISTERS_35_19_port, REGISTERS_35_18_port, 
      REGISTERS_35_17_port, REGISTERS_35_16_port, REGISTERS_35_15_port, 
      REGISTERS_35_14_port, REGISTERS_35_13_port, REGISTERS_35_12_port, 
      REGISTERS_35_11_port, REGISTERS_35_10_port, REGISTERS_35_9_port, 
      REGISTERS_35_8_port, REGISTERS_35_7_port, REGISTERS_35_6_port, 
      REGISTERS_35_5_port, REGISTERS_35_4_port, REGISTERS_35_3_port, 
      REGISTERS_35_2_port, REGISTERS_35_1_port, REGISTERS_35_0_port, 
      REGISTERS_36_31_port, REGISTERS_36_30_port, REGISTERS_36_29_port, 
      REGISTERS_36_28_port, REGISTERS_36_27_port, REGISTERS_36_26_port, 
      REGISTERS_36_25_port, REGISTERS_36_24_port, REGISTERS_36_23_port, 
      REGISTERS_36_22_port, REGISTERS_36_21_port, REGISTERS_36_20_port, 
      REGISTERS_36_19_port, REGISTERS_36_18_port, REGISTERS_36_17_port, 
      REGISTERS_36_16_port, REGISTERS_36_15_port, REGISTERS_36_14_port, 
      REGISTERS_36_13_port, REGISTERS_36_12_port, REGISTERS_36_11_port, 
      REGISTERS_36_10_port, REGISTERS_36_9_port, REGISTERS_36_8_port, 
      REGISTERS_36_7_port, REGISTERS_36_6_port, REGISTERS_36_5_port, 
      REGISTERS_36_4_port, REGISTERS_36_3_port, REGISTERS_36_2_port, 
      REGISTERS_36_1_port, REGISTERS_36_0_port, REGISTERS_37_31_port, 
      REGISTERS_37_30_port, REGISTERS_37_29_port, REGISTERS_37_28_port, 
      REGISTERS_37_27_port, REGISTERS_37_26_port, REGISTERS_37_25_port, 
      REGISTERS_37_24_port, REGISTERS_37_23_port, REGISTERS_37_22_port, 
      REGISTERS_37_21_port, REGISTERS_37_20_port, REGISTERS_37_19_port, 
      REGISTERS_37_18_port, REGISTERS_37_17_port, REGISTERS_37_16_port, 
      REGISTERS_37_15_port, REGISTERS_37_14_port, REGISTERS_37_13_port, 
      REGISTERS_37_12_port, REGISTERS_37_11_port, REGISTERS_37_10_port, 
      REGISTERS_37_9_port, REGISTERS_37_8_port, REGISTERS_37_7_port, 
      REGISTERS_37_6_port, REGISTERS_37_5_port, REGISTERS_37_4_port, 
      REGISTERS_37_3_port, REGISTERS_37_2_port, REGISTERS_37_1_port, 
      REGISTERS_37_0_port, REGISTERS_38_31_port, REGISTERS_38_30_port, 
      REGISTERS_38_29_port, REGISTERS_38_28_port, REGISTERS_38_27_port, 
      REGISTERS_38_26_port, REGISTERS_38_25_port, REGISTERS_38_24_port, 
      REGISTERS_38_23_port, REGISTERS_38_22_port, REGISTERS_38_21_port, 
      REGISTERS_38_20_port, REGISTERS_38_19_port, REGISTERS_38_18_port, 
      REGISTERS_38_17_port, REGISTERS_38_16_port, REGISTERS_38_15_port, 
      REGISTERS_38_14_port, REGISTERS_38_13_port, REGISTERS_38_12_port, 
      REGISTERS_38_11_port, REGISTERS_38_10_port, REGISTERS_38_9_port, 
      REGISTERS_38_8_port, REGISTERS_38_7_port, REGISTERS_38_6_port, 
      REGISTERS_38_5_port, REGISTERS_38_4_port, REGISTERS_38_3_port, 
      REGISTERS_38_2_port, REGISTERS_38_1_port, REGISTERS_38_0_port, 
      REGISTERS_39_31_port, REGISTERS_39_30_port, REGISTERS_39_29_port, 
      REGISTERS_39_28_port, REGISTERS_39_27_port, REGISTERS_39_26_port, 
      REGISTERS_39_25_port, REGISTERS_39_24_port, REGISTERS_39_23_port, 
      REGISTERS_39_22_port, REGISTERS_39_21_port, REGISTERS_39_20_port, 
      REGISTERS_39_19_port, REGISTERS_39_18_port, REGISTERS_39_17_port, 
      REGISTERS_39_16_port, REGISTERS_39_15_port, REGISTERS_39_14_port, 
      REGISTERS_39_13_port, REGISTERS_39_12_port, REGISTERS_39_11_port, 
      REGISTERS_39_10_port, REGISTERS_39_9_port, REGISTERS_39_8_port, 
      REGISTERS_39_7_port, REGISTERS_39_6_port, REGISTERS_39_5_port, 
      REGISTERS_39_4_port, REGISTERS_39_3_port, REGISTERS_39_2_port, 
      REGISTERS_39_1_port, REGISTERS_39_0_port, N4389, N4390, N4391, N4392, 
      N4393, N4394, N4395, N4396, N4397, N4398, N4399, N4400, N4401, N4402, 
      N4403, N4404, N4405, N4406, N4407, N4408, N4409, N4410, N4411, N4412, 
      N4413, N4414, N4415, N4416, N4417, N4418, N4419, N4420, N4495, N4496, 
      N4497, N4498, N4499, N4500, N4501, N4502, N4503, N4504, N4505, N4506, 
      N4507, N4508, N4509, N4510, N4511, N4512, N4513, N4514, N4515, N4516, 
      N4517, N4518, N4519, N4520, N4521, N4522, N4523, N4524, N4525, N4526, 
      SWP_31_port, SWP_30_port, SWP_29_port, SWP_28_port, SWP_27_port, 
      SWP_26_port, SWP_25_port, SWP_24_port, SWP_23_port, SWP_22_port, 
      SWP_21_port, SWP_20_port, SWP_19_port, SWP_18_port, SWP_17_port, 
      SWP_16_port, SWP_15_port, SWP_14_port, SWP_13_port, SWP_12_port, 
      SWP_11_port, SWP_10_port, SWP_9_port, SWP_8_port, SWP_7_port, SWP_6_port,
      SWP_5_port, SWP_4_port, SWP_3_port, SWP_1_port, SWP_0_port, N5250, N5251,
      N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, 
      N5262, N5263, N5264, N5265, N5266, N5267, N5268, N5269, N5270, N5271, 
      N5272, N5273, N5274, N5275, N5276, N5277, N5278, N5279, N5280, N5281, 
      N12205, N12206, N12207, N12208, N12209, N12210, N12211, N12212, N12213, 
      N12214, N12215, N12216, N12217, N12218, N12219, N12220, N12221, N12222, 
      N12223, N12224, N12225, N12226, N12227, N12228, N12229, N12230, N12231, 
      N12232, N12233, N12234, N12235, N12236, N12237, N12238, N12239, N12240, 
      N12241, N12242, N12243, N12244, N12245, N12246, N12247, N12248, N12249, 
      N12250, N12251, N12252, N12253, N12254, N12255, N12256, N12257, N12258, 
      N12259, N12260, N12261, N12262, N12263, N12264, N12265, N12266, N12267, 
      N12268, N12269, N12270, N12271, N12272, N12273, N12274, N12275, N12276, 
      N12277, N12278, N12279, N12280, N12281, N12282, N12283, N12284, N12285, 
      N12286, N12287, N12288, N12289, N12290, N12291, N12292, N12293, N12294, 
      N12295, N12296, N12297, N12298, N12299, N12300, N13831, N13832, N13833, 
      N13834, N13835, N13836, N13837, N13838, N13839, N13840, N13841, N13842, 
      N13843, N13844, N13845, N13846, N13847, N13848, N13849, N13850, N13851, 
      N13852, N13853, N13854, N13855, N13856, N13857, N13858, N13859, N13860, 
      N13861, N13862, N50337, N50338, N50340, N50341, N50342, N50343, N50344, 
      N50345, N50346, N50347, N50348, N50349, N50350, N50351, N50352, N50353, 
      N50354, N50355, N50356, N50357, N50358, N50359, N50360, N50361, N50362, 
      N50363, N50364, N50365, N50366, N50367, N50368, n49, n52, n55, n58, n61, 
      n62, n65, n89, n90, n10323, n10324, n10325, n10326, n10327, n10328, 
      n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, 
      n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, 
      n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, 
      n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, 
      n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, 
      n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, 
      n10383, n10384, n10385, n10386, n10388, n10389, n10390, n10391, n10392, 
      n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, 
      n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, 
      n10411, n10412, n10413, n10446, n10447, n10448, n10449, n10450, n10451, 
      n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, 
      n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, 
      n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, 
      n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, 
      n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, 
      n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, 
      n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, 
      n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, 
      n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, 
      n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, 
      n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, 
      n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, 
      n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, 
      n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, 
      n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, 
      n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, 
      n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, 
      n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, 
      n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, 
      n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, 
      n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, 
      n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, 
      n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, 
      n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, 
      n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, 
      n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, 
      n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, 
      n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, 
      n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, 
      n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, 
      n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, 
      n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, 
      n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, 
      n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, 
      n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, 
      n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, 
      n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, 
      n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, 
      n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, 
      n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, 
      n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, 
      n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, 
      n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, 
      n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, 
      n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, 
      n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, 
      n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, 
      n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, 
      n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, 
      n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, 
      n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, 
      n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, 
      n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, 
      n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, 
      n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, 
      n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, 
      n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, 
      n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, 
      n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, 
      n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, 
      n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, 
      n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, 
      n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, 
      n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, 
      n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, 
      n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, 
      n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, 
      n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, 
      n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, 
      n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, 
      n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, 
      n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, 
      n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, 
      n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, 
      n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, 
      n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, 
      n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, 
      n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, 
      n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, 
      n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, 
      n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, 
      n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, 
      n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, 
      n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, 
      n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, 
      n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, 
      n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, 
      n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, 
      n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, 
      n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, 
      n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, 
      n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, 
      n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, 
      n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, 
      n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, 
      n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, 
      n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, 
      n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
      n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, 
      n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, 
      n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, 
      n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, 
      n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, 
      n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, 
      n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, 
      n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, 
      n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, 
      n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, 
      n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, 
      n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, 
      n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, 
      n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, 
      n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, 
      n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, 
      n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, 
      n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, 
      n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, 
      n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, 
      n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, 
      n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, 
      n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, 
      n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, 
      n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, 
      n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, 
      n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, 
      n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, 
      n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, 
      n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, 
      n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, 
      n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, 
      n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, 
      n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, 
      n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, 
      n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, 
      n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, 
      n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, 
      n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, 
      n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, 
      n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, 
      n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, 
      n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, 
      n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, 
      n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, 
      n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, 
      n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, 
      n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, 
      n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, 
      n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, 
      n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, 
      n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, 
      n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, 
      n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, 
      n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, 
      n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, 
      n11838, n11839, n11840, n11841, n11842, n11859, n11860, n11861, n11862, 
      n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11872, n11873, 
      n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, 
      n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, 
      n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, 
      n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, 
      n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, 
      n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, 
      n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, 
      n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, 
      n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, 
      n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, 
      n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, 
      n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, 
      n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, 
      n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, 
      n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, 
      n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, 
      n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, 
      n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, 
      n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, 
      n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, 
      n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, 
      n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, 
      n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, 
      n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, 
      n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, 
      n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, 
      n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, 
      n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, 
      n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, 
      n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, 
      n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, 
      n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, 
      n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, 
      n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, 
      n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, 
      n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, 
      n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205_port, 
      n12206_port, n12207_port, n12208_port, n12209_port, n12210_port, 
      n12211_port, n12212_port, n12213_port, n12214_port, n12215_port, 
      n12216_port, n12217_port, n12218_port, n12219_port, n12220_port, 
      n12221_port, n12222_port, n12223_port, n12224_port, n12225_port, 
      n12226_port, n12227_port, n12228_port, n12229_port, n12230_port, 
      n12231_port, n12232_port, n12233_port, n12234_port, n12235_port, 
      n12236_port, n12237_port, n12238_port, n12239_port, n12240_port, 
      n12241_port, n12242_port, n12243_port, n12244_port, n12245_port, 
      n12246_port, n12247_port, n12248_port, n12249_port, n12250_port, 
      n12251_port, n12252_port, n12253_port, n12254_port, n12255_port, 
      n12256_port, n12257_port, n12258_port, n12259_port, n12260_port, 
      n12261_port, n12262_port, n12263_port, n12264_port, n12265_port, 
      n12266_port, n12267_port, n12268_port, n12269_port, n12270_port, 
      n12271_port, n12272_port, n12273_port, n12274_port, n12275_port, 
      n12276_port, n12277_port, n12278_port, n12279_port, n12280_port, 
      n12281_port, n12282_port, n12283_port, n12284_port, n12285_port, 
      n12286_port, n12287_port, n12288_port, n12289_port, n12290_port, 
      n12291_port, n12292_port, n12293_port, n12294_port, n12295_port, 
      n12296_port, n12297_port, n12298_port, n12299_port, n12300_port, n12301, 
      n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, 
      n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, 
      n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, 
      n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, 
      n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, 
      n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, 
      n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, 
      n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, 
      n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, 
      n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, 
      n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, 
      n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, 
      n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, 
      n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, 
      n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, 
      n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, 
      n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, 
      n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, 
      n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, 
      n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, 
      n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, 
      n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, 
      n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, 
      n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, 
      n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, 
      n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, 
      n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, 
      n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, 
      n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, 
      n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, 
      n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, 
      n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, 
      n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, 
      n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, 
      n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, 
      n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, 
      n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, 
      n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, 
      n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, 
      n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, 
      n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, 
      n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, 
      n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, 
      n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, 
      n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, 
      n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, 
      n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, 
      n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, 
      n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, 
      n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, 
      n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, 
      n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, 
      n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, 
      n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, 
      n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, 
      n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, 
      n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, 
      n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, 
      n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, 
      n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, 
      n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, 
      n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, 
      n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, 
      n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, 
      n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, 
      n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, 
      n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, 
      n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, 
      n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, 
      n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, 
      n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, 
      n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, 
      n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, 
      n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, 
      n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, 
      n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, 
      n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, 
      n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, 
      n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, 
      n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, 
      n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, 
      n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, 
      n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, 
      n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, 
      n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, 
      n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, 
      n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, 
      n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, 
      n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, 
      n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, 
      n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, 
      n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, 
      n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, 
      n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, 
      n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, 
      n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, 
      n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, 
      n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, 
      n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, 
      r3007_A_0_port, r3007_A_1_port, r3007_A_2_port, r3007_A_3_port, 
      r3007_A_4_port, r3013_A_0_port, r3013_A_1_port, r3013_A_2_port, 
      r3013_A_3_port, r3013_A_4_port, sub_65_carry_4_port, sub_64_carry_4_port,
      sub_63_carry_4_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60
      , n63, n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
      n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
      n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
      n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
      n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
      n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
      n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
      n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564_port, n3565_port, 
      n3566_port, n3567_port, n3568_port, n3569_port, n3570_port, n3571_port, 
      n3572_port, n3573, n3574, n3575, n3576, n3577_port, n3578_port, 
      n3579_port, n3580_port, n3581_port, n3582_port, n3583_port, n3584_port, 
      n3585_port, n3586, n3587, n3588, n3589, n3590_port, n3591_port, 
      n3592_port, n3593_port, n3594_port, n3595_port, n3596_port, n3597_port, 
      n3598_port, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607
      , n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, 
      n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, 
      n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, 
      n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, 
      n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, 
      n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, 
      n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, 
      n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, 
      n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, 
      n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, 
      n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, 
      n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, 
      n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, 
      n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, 
      n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, 
      n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, 
      n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, 
      n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, 
      n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, 
      n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, 
      n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, 
      n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, 
      n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, 
      n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, 
      n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, 
      n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, 
      n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, 
      n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, 
      n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, 
      n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, 
      n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, 
      n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, 
      n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, 
      n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, 
      n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, 
      n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, 
      n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, 
      n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, 
      n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, 
      n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, 
      n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, 
      n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, 
      n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
      n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
      n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
      n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
      n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, 
      n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
      n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, 
      n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, 
      n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, 
      n4388, n4389_port, n4390_port, n4391_port, n4392_port, n4393_port, 
      n4394_port, n4395_port, n4396_port, n4397_port, n4398_port, n4399_port, 
      n4400_port, n4401_port, n4402_port, n4403_port, n4404_port, n4405_port, 
      n4406_port, n4407_port, n4408_port, n4409_port, n4410_port, n4411_port, 
      n4412_port, n4413_port, n4414_port, n4415_port, n4416_port, n4417_port, 
      n4418_port, n4419_port, n4420_port, n4421, n4422, n4423, n4424, n4425, 
      n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, 
      n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, 
      n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, 
      n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, 
      n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, 
      n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, 
      n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495_port
      , n4496_port, n4497_port, n4498_port, n4499_port, n4500_port, n4501_port,
      n4502_port, n4503_port, n4504_port, n4505_port, n4506_port, n4507_port, 
      n4508_port, n4509_port, n4510_port, n4511_port, n4512_port, n4513_port, 
      n4514_port, n4515_port, n4516_port, n4517_port, n4518_port, n4519_port, 
      n4520_port, n4521_port, n4522_port, n4523_port, n4524_port, n4525_port, 
      n4526_port, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535
      , n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, 
      n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, 
      n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, 
      n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, 
      n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, 
      n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, 
      n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, 
      n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, 
      n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, 
      n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, 
      n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, 
      n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, 
      n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, 
      n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, 
      n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, 
      n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, 
      n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, 
      n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, 
      n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, 
      n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, 
      n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, 
      n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, 
      n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, 
      n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, 
      n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, 
      n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, 
      n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, 
      n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, 
      n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, 
      n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, 
      n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, 
      n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, 
      n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, 
      n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, 
      n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, 
      n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, 
      n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, 
      n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, 
      n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, 
      n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, 
      n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, 
      n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, 
      n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, 
      n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, 
      n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, 
      n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, 
      n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, 
      n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, 
      n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, 
      n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, 
      n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, 
      n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, 
      n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, 
      n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, 
      n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, 
      n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, 
      n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, 
      n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, 
      n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
      n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, 
      n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, 
      n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, 
      n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, 
      n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, 
      n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, 
      n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, 
      n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, 
      n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, 
      n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, 
      n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, 
      n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, 
      n5246, n5247, n5248, n5249, n5250_port, n5251_port, n5252_port, 
      n5253_port, n5254_port, n5255_port, n5256_port, n5257_port, n5258_port, 
      n5259_port, n5260_port, n5261_port, n5262_port, n5263_port, n5264_port, 
      n5265_port, n5266_port, n5267_port, n5268_port, n5269_port, n5270_port, 
      n5271_port, n5272_port, n5273_port, n5274_port, n5275_port, n5276_port, 
      n5277_port, n5278_port, n5279_port, n5280_port, n5281_port, n5282, n5283,
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, 
      n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, 
      n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, 
      n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, 
      n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, 
      n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, 
      n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, 
      n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, 
      n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, 
      n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, 
      n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, 
      n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
      n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, 
      n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, 
      n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, 
      n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, 
      n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, 
      n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, 
      n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, 
      n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, 
      n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, 
      n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, 
      n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, 
      n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
      n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, 
      n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, 
      n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, 
      n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, 
      n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, 
      n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, 
      n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, 
      n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, 
      n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, 
      n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, 
      n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, 
      n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, 
      n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, 
      n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, 
      n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, 
      n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, 
      n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, 
      n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, 
      n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, 
      n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, 
      n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, 
      n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, 
      n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, 
      n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, 
      n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, 
      n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, 
      n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, 
      n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, 
      n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, 
      n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, 
      n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
      n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, 
      n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, 
      n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, 
      n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
      n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
      n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, 
      n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, 
      n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, 
      n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
      n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, 
      n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, 
      n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, 
      n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, 
      n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, 
      n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, 
      n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, 
      n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, 
      n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, 
      n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
      n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, 
      n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, 
      n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, 
      n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, 
      n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, 
      n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, 
      n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, 
      n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, 
      n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, 
      n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, 
      n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, 
      n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
      n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, 
      n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, 
      n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, 
      n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
      n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, 
      n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, 
      n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, 
      n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, 
      n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, 
      n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, 
      n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
      n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, 
      n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
      n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, 
      n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, 
      n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, 
      n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, 
      n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, 
      n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, 
      n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
      n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, 
      n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
      n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
      n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
      n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, 
      n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, 
      n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
      n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, 
      n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, 
      n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, 
      n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
      n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, 
      n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, 
      n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
      n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, 
      n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
      n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, 
      n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
      n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, 
      n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, 
      n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
      n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
      n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, 
      n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, 
      n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
      n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, 
      n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, 
      n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, 
      n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
      n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, 
      n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, 
      n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, 
      n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, 
      n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, 
      n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, 
      n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, 
      n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, 
      n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
      n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, 
      n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
      n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, 
      n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
      n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, 
      n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
      n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
      n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, 
      n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, 
      n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
      n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, 
      n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, 
      n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
      n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, 
      n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, 
      n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, 
      n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, 
      n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, 
      n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, 
      n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, 
      n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, 
      n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, 
      n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, 
      n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, 
      n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, 
      n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, 
      n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, 
      n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, 
      n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, 
      n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, 
      n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
      n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
      n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, 
      n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, 
      n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
      n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, 
      n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
      n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, 
      n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, 
      n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, 
      n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
      n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, 
      n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
      n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, 
      n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, 
      n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, 
      n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, 
      n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, 
      n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, 
      n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, 
      n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, 
      n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, 
      n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, 
      n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, 
      n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, 
      n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, 
      n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, 
      n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, 
      n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, 
      n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, 
      n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, 
      n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, 
      n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
      n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, 
      n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, 
      n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, 
      n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, 
      n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, 
      n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, 
      n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, 
      n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, 
      n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, 
      n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, 
      n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, 
      n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, 
      n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, 
      n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, 
      n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, 
      n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, 
      n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, 
      n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, 
      n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, 
      n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, 
      n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, 
      n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, 
      n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, 
      n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, 
      n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, 
      n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, 
      n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, 
      n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, 
      n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
      n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, 
      n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, 
      n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, 
      n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, 
      n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, 
      n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, 
      n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, 
      n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, 
      n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, 
      n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, 
      n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, 
      n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, 
      n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, 
      n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, 
      n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, 
      n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, 
      n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, 
      n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
      n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, 
      n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, 
      n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, 
      n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, 
      n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, 
      n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, 
      n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, 
      n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, 
      n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, 
      n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, 
      n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, 
      n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, 
      n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, 
      n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, 
      n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, 
      n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, 
      n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, 
      n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, 
      n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, 
      n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, 
      n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, 
      n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, 
      n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, 
      n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, 
      n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, 
      n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, 
      n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, 
      n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, 
      n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, 
      n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, 
      n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, 
      n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, 
      n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, 
      n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, 
      n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, 
      n10319, n10320, n10321, n10322, n10387, n10414, n10415, n10416, n10417, 
      n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, 
      n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, 
      n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, 
      n10445, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, 
      n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11870, 
      n11871, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, 
      n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, 
      n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, 
      n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, 
      n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, 
      n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, 
      n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, 
      n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, 
      n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, 
      n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, 
      n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, 
      n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, 
      n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, 
      n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, 
      n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, 
      n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, 
      n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, 
      n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, 
      n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, 
      n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, 
      n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, 
      n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, 
      n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, 
      n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, 
      n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, 
      n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, 
      n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, 
      n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, 
      n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, 
      n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, 
      n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, 
      n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, 
      n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, 
      n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, 
      n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, 
      n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, 
      n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, 
      n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, 
      n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, 
      n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, 
      n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, 
      n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, 
      n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, 
      n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, 
      n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, 
      n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, 
      n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, 
      n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, 
      n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, 
      n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, 
      n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, 
      n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, 
      n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, 
      n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, 
      n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, 
      n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, 
      n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, 
      n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, 
      n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, 
      n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, 
      n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, 
      n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, 
      n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, 
      n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, 
      n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, 
      n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, 
      n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, 
      n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, 
      n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, 
      n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, 
      n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, 
      n13831_port, n13832_port, n13833_port, n13834_port, n13835_port, 
      n13836_port, n13837_port, n13838_port, n13839_port, n13840_port, 
      n13841_port, n13842_port, n13843_port, n13844_port, n13845_port, 
      n13846_port, n13847_port, n13848_port, n13849_port, n13850_port, 
      n13851_port, n13852_port, n13853_port, n13854_port, n13855_port, 
      n13856_port, n13857_port, n13858_port, n13859_port, n13860_port, 
      n13861_port, n13862_port, n13863, n13864, n13865, n13866, n13867, n13868,
      n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, 
      n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, 
      n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, 
      n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, 
      n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, 
      n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, 
      n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, 
      n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, 
      n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, 
      n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, 
      n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, 
      n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, 
      n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, 
      n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, 
      n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, 
      n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, 
      n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, 
      n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, 
      n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, 
      n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, 
      n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, 
      n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, 
      n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, 
      n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, 
      n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, 
      n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, 
      n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, 
      n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, 
      n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, 
      n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, 
      n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, 
      n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, 
      n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, 
      n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, 
      n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, 
      n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, 
      n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, 
      n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, 
      n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, 
      n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, 
      n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, 
      n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, 
      n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, 
      n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, 
      n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, 
      n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, 
      n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, 
      n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, 
      n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, 
      n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, 
      n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, 
      n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, 
      n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, 
      n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, 
      n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, 
      n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, 
      n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, 
      n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, 
      n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, 
      n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, 
      n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, 
      n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, 
      n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, 
      n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, 
      n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, 
      n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, 
      n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, 
      n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, 
      n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, 
      n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, 
      n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, 
      n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, 
      n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, 
      n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, 
      n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, 
      n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, 
      n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, 
      n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, 
      n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, 
      n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, 
      n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, 
      n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, 
      n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, 
      n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, 
      n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, 
      n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, 
      n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, 
      n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, 
      n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, 
      n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, 
      n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, 
      n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, 
      n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, 
      n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, 
      n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, 
      n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, 
      n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, 
      n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, 
      n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, 
      n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, 
      n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, 
      n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, 
      n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, 
      n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, 
      n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, 
      n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, 
      n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, 
      n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, 
      n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, 
      n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, 
      n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, 
      n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, 
      n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, 
      n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, 
      n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, 
      n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, 
      n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, 
      n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, 
      n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, 
      n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, 
      n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, 
      n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, 
      n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, 
      n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, 
      n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, 
      n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, 
      n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, 
      n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, 
      n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, 
      n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, 
      n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, 
      n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, 
      n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, 
      n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, 
      n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, 
      n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, 
      n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, 
      n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, 
      n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, 
      n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, 
      n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, 
      n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, 
      n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, 
      n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, 
      n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, 
      n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, 
      n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, 
      n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, 
      n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, 
      n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, 
      n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, 
      n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, 
      n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, 
      n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, 
      n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, 
      n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, 
      n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, 
      n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, 
      n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, 
      n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, 
      n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, 
      n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, 
      n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, 
      n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, 
      n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, 
      n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, 
      n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, 
      n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, 
      n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, 
      n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, 
      n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, 
      n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, 
      n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, 
      n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, 
      n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, 
      n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, 
      n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, 
      n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, 
      n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, 
      n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, 
      n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, 
      n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, 
      n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, 
      n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, 
      n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, 
      n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, 
      n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, 
      n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, 
      n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, 
      n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, 
      n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, 
      n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, 
      n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, 
      n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, 
      n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, 
      n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, 
      n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, 
      n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, 
      n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, 
      n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, 
      n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, 
      n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, 
      n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, 
      n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, 
      n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, 
      n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, 
      n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, 
      n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, 
      n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, 
      n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, 
      n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, 
      n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, 
      n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, 
      n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, 
      n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, 
      n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, 
      n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, 
      n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, 
      n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, 
      n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, 
      n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, 
      n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, 
      n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, 
      n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, 
      n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, 
      n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, 
      n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, 
      n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, 
      n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, 
      n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, 
      n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, 
      n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, 
      n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, 
      n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, 
      n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, 
      n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, 
      n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, 
      n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, 
      n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, 
      n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, 
      n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, 
      n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, 
      n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, 
      n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, 
      n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, 
      n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, 
      n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, 
      n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, 
      n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, 
      n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, 
      n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, 
      n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, 
      n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, 
      n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, 
      n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, 
      n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, 
      n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, 
      n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, 
      n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, 
      n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, 
      n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, 
      n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, 
      n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, 
      n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, 
      n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, 
      n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, 
      n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, 
      n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, 
      n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, 
      n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, 
      n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, 
      n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, 
      n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, 
      n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, 
      n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, 
      n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, 
      n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, 
      n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, 
      n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, 
      n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, 
      n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, 
      n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, 
      n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, 
      n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, 
      n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, 
      n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, 
      n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, 
      n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, 
      n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, 
      n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, 
      n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510 : std_logic;

begin
   FILL <= FILL_port;
   MEM_OUT <= ( MEM_OUT_31_port, MEM_OUT_30_port, MEM_OUT_29_port, 
      MEM_OUT_28_port, MEM_OUT_27_port, MEM_OUT_26_port, MEM_OUT_25_port, 
      MEM_OUT_24_port, MEM_OUT_23_port, MEM_OUT_22_port, MEM_OUT_21_port, 
      MEM_OUT_20_port, MEM_OUT_19_port, MEM_OUT_18_port, MEM_OUT_17_port, 
      MEM_OUT_16_port, MEM_OUT_15_port, MEM_OUT_14_port, MEM_OUT_13_port, 
      MEM_OUT_12_port, MEM_OUT_11_port, MEM_OUT_10_port, MEM_OUT_9_port, 
      MEM_OUT_8_port, MEM_OUT_7_port, MEM_OUT_6_port, MEM_OUT_5_port, 
      MEM_OUT_4_port, MEM_OUT_3_port, MEM_OUT_2_port, MEM_OUT_1_port, 
      MEM_OUT_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n49 <= '0';
   n52 <= '0';
   n55 <= '0';
   n58 <= '0';
   n61 <= '0';
   n62 <= '0';
   n65 <= '0';
   fspill_reg : DFF_X1 port map( D => n13192, CK => n978, Q => n16455, QN => 
                           n116);
   canrestore_reg_0_inst : DFF_X1 port map( D => n13159, CK => n978, Q => n117,
                           QN => n_1469);
   CWP_reg_31_inst : DFF_X1 port map( D => n13191, CK => n977, Q => CWP_31_port
                           , QN => n11790);
   CWP_reg_2_inst : DFF_X1 port map( D => n13188, CK => n978, Q => CWP_2_port, 
                           QN => n11861);
   CWP_reg_30_inst : DFF_X1 port map( D => n13160, CK => n972, Q => CWP_30_port
                           , QN => n11817);
   CWP_reg_3_inst : DFF_X1 port map( D => n13187, CK => n977, Q => CWP_3_port, 
                           QN => n11860);
   CWP_reg_29_inst : DFF_X1 port map( D => n13161, CK => n972, Q => CWP_29_port
                           , QN => n11818);
   CWP_reg_4_inst : DFF_X1 port map( D => n13186, CK => n977, Q => CWP_4_port, 
                           QN => n11859);
   CWP_reg_28_inst : DFF_X1 port map( D => n13162, CK => n972, Q => CWP_28_port
                           , QN => n11819);
   CWP_reg_27_inst : DFF_X1 port map( D => n13163, CK => n972, Q => CWP_27_port
                           , QN => n11820);
   CWP_reg_26_inst : DFF_X1 port map( D => n13164, CK => n972, Q => CWP_26_port
                           , QN => n11821);
   CWP_reg_25_inst : DFF_X1 port map( D => n13165, CK => n972, Q => CWP_25_port
                           , QN => n11822);
   CWP_reg_24_inst : DFF_X1 port map( D => n13166, CK => n972, Q => CWP_24_port
                           , QN => n11823);
   CWP_reg_23_inst : DFF_X1 port map( D => n13167, CK => n973, Q => CWP_23_port
                           , QN => n11824);
   CWP_reg_22_inst : DFF_X1 port map( D => n13168, CK => n973, Q => CWP_22_port
                           , QN => n11825);
   CWP_reg_21_inst : DFF_X1 port map( D => n13169, CK => n973, Q => CWP_21_port
                           , QN => n11826);
   CWP_reg_20_inst : DFF_X1 port map( D => n13170, CK => n973, Q => CWP_20_port
                           , QN => n11827);
   CWP_reg_19_inst : DFF_X1 port map( D => n13171, CK => n973, Q => CWP_19_port
                           , QN => n11828);
   CWP_reg_18_inst : DFF_X1 port map( D => n13172, CK => n973, Q => CWP_18_port
                           , QN => n11829);
   CWP_reg_17_inst : DFF_X1 port map( D => n13173, CK => n973, Q => CWP_17_port
                           , QN => n11830);
   CWP_reg_16_inst : DFF_X1 port map( D => n13174, CK => n973, Q => CWP_16_port
                           , QN => n11831);
   CWP_reg_15_inst : DFF_X1 port map( D => n13175, CK => n973, Q => CWP_15_port
                           , QN => n11832);
   CWP_reg_14_inst : DFF_X1 port map( D => n13176, CK => n973, Q => CWP_14_port
                           , QN => n11833);
   CWP_reg_13_inst : DFF_X1 port map( D => n13177, CK => n973, Q => CWP_13_port
                           , QN => n11834);
   CWP_reg_12_inst : DFF_X1 port map( D => n13178, CK => n974, Q => CWP_12_port
                           , QN => n11835);
   CWP_reg_11_inst : DFF_X1 port map( D => n13179, CK => n974, Q => CWP_11_port
                           , QN => n11836);
   CWP_reg_10_inst : DFF_X1 port map( D => n13180, CK => n974, Q => CWP_10_port
                           , QN => n11837);
   CWP_reg_9_inst : DFF_X1 port map( D => n13181, CK => n974, Q => CWP_9_port, 
                           QN => n11838);
   CWP_reg_8_inst : DFF_X1 port map( D => n13182, CK => n974, Q => CWP_8_port, 
                           QN => n11839);
   CWP_reg_7_inst : DFF_X1 port map( D => n13183, CK => n974, Q => CWP_7_port, 
                           QN => n11840);
   CWP_reg_6_inst : DFF_X1 port map( D => n13184, CK => n974, Q => CWP_6_port, 
                           QN => n11841);
   CWP_reg_5_inst : DFF_X1 port map( D => n13185, CK => n974, Q => CWP_5_port, 
                           QN => n11842);
   CWP_reg_1_inst : DFF_X1 port map( D => n13189, CK => n972, Q => CWP_1_port, 
                           QN => n11862);
   CWP_reg_0_inst : DFF_X1 port map( D => n13190, CK => n972, Q => CWP_0_port, 
                           QN => n11863);
   SWP_reg_0_inst : DFF_X1 port map( D => n13158, CK => n974, Q => SWP_0_port, 
                           QN => n11869);
   SWP_reg_31_inst : DFF_X1 port map( D => n11816, CK => n975, Q => SWP_31_port
                           , QN => n10413);
   SWP_reg_1_inst : DFF_X1 port map( D => n13157, CK => n974, Q => SWP_1_port, 
                           QN => n11868);
   SWP_reg_2_inst : DFF_X1 port map( D => n13156, CK => n977, Q => n1, QN => 
                           n11867);
   SWP_reg_4_inst : DFF_X1 port map( D => n13154, CK => n977, Q => SWP_4_port, 
                           QN => n11865);
   SWP_reg_5_inst : DFF_X1 port map( D => n13153, CK => n977, Q => SWP_5_port, 
                           QN => n11864);
   SWP_reg_6_inst : DFF_X1 port map( D => n11791, CK => n977, Q => SWP_6_port, 
                           QN => n10388);
   SWP_reg_7_inst : DFF_X1 port map( D => n11792, CK => n977, Q => SWP_7_port, 
                           QN => n10389);
   SWP_reg_8_inst : DFF_X1 port map( D => n11793, CK => n977, Q => SWP_8_port, 
                           QN => n10390);
   SWP_reg_9_inst : DFF_X1 port map( D => n11794, CK => n977, Q => SWP_9_port, 
                           QN => n10391);
   SWP_reg_10_inst : DFF_X1 port map( D => n11795, CK => n976, Q => SWP_10_port
                           , QN => n10392);
   SWP_reg_11_inst : DFF_X1 port map( D => n11796, CK => n976, Q => SWP_11_port
                           , QN => n10393);
   SWP_reg_12_inst : DFF_X1 port map( D => n11797, CK => n976, Q => SWP_12_port
                           , QN => n10394);
   SWP_reg_13_inst : DFF_X1 port map( D => n11798, CK => n976, Q => SWP_13_port
                           , QN => n10395);
   SWP_reg_14_inst : DFF_X1 port map( D => n11799, CK => n976, Q => SWP_14_port
                           , QN => n10396);
   SWP_reg_15_inst : DFF_X1 port map( D => n11800, CK => n976, Q => SWP_15_port
                           , QN => n10397);
   SWP_reg_16_inst : DFF_X1 port map( D => n11801, CK => n976, Q => SWP_16_port
                           , QN => n10398);
   SWP_reg_17_inst : DFF_X1 port map( D => n11802, CK => n976, Q => SWP_17_port
                           , QN => n10399);
   SWP_reg_18_inst : DFF_X1 port map( D => n11803, CK => n976, Q => SWP_18_port
                           , QN => n10400);
   SWP_reg_19_inst : DFF_X1 port map( D => n11804, CK => n976, Q => SWP_19_port
                           , QN => n10401);
   SWP_reg_20_inst : DFF_X1 port map( D => n11805, CK => n976, Q => SWP_20_port
                           , QN => n10402);
   SWP_reg_21_inst : DFF_X1 port map( D => n11806, CK => n975, Q => SWP_21_port
                           , QN => n10403);
   SWP_reg_22_inst : DFF_X1 port map( D => n11807, CK => n975, Q => SWP_22_port
                           , QN => n10404);
   SWP_reg_23_inst : DFF_X1 port map( D => n11808, CK => n975, Q => SWP_23_port
                           , QN => n10405);
   SWP_reg_24_inst : DFF_X1 port map( D => n11809, CK => n975, Q => SWP_24_port
                           , QN => n10406);
   SWP_reg_25_inst : DFF_X1 port map( D => n11810, CK => n975, Q => SWP_25_port
                           , QN => n10407);
   SWP_reg_26_inst : DFF_X1 port map( D => n11811, CK => n975, Q => SWP_26_port
                           , QN => n10408);
   SWP_reg_27_inst : DFF_X1 port map( D => n11812, CK => n975, Q => SWP_27_port
                           , QN => n10409);
   SWP_reg_28_inst : DFF_X1 port map( D => n11813, CK => n975, Q => SWP_28_port
                           , QN => n10410);
   SWP_reg_29_inst : DFF_X1 port map( D => n11814, CK => n975, Q => SWP_29_port
                           , QN => n10411);
   SWP_reg_30_inst : DFF_X1 port map( D => n11815, CK => n975, Q => SWP_30_port
                           , QN => n10412);
   OUT2_reg_31_inst : DFF_X1 port map( D => n10447, CK => n953, Q => OUT2(31), 
                           QN => n10386);
   OUT2_reg_30_inst : DFF_X1 port map( D => n10450, CK => n895, Q => OUT2(30), 
                           QN => n10385);
   OUT2_reg_29_inst : DFF_X1 port map( D => n10453, CK => n892, Q => OUT2(29), 
                           QN => n10384);
   OUT2_reg_28_inst : DFF_X1 port map( D => n10456, CK => n957, Q => OUT2(28), 
                           QN => n10383);
   OUT2_reg_27_inst : DFF_X1 port map( D => n10459, CK => n937, Q => OUT2(27), 
                           QN => n10382);
   OUT2_reg_26_inst : DFF_X1 port map( D => n10462, CK => n934, Q => OUT2(26), 
                           QN => n10381);
   OUT2_reg_25_inst : DFF_X1 port map( D => n10465, CK => n930, Q => OUT2(25), 
                           QN => n10380);
   OUT2_reg_24_inst : DFF_X1 port map( D => n10468, CK => n941, Q => OUT2(24), 
                           QN => n10379);
   OUT2_reg_23_inst : DFF_X1 port map( D => n10471, CK => n926, Q => OUT2(23), 
                           QN => n10378);
   OUT2_reg_22_inst : DFF_X1 port map( D => n10474, CK => n922, Q => OUT2(22), 
                           QN => n10377);
   OUT2_reg_21_inst : DFF_X1 port map( D => n10477, CK => n918, Q => OUT2(21), 
                           QN => n10376);
   OUT2_reg_20_inst : DFF_X1 port map( D => n10480, CK => n915, Q => OUT2(20), 
                           QN => n10375);
   OUT2_reg_19_inst : DFF_X1 port map( D => n10483, CK => n911, Q => OUT2(19), 
                           QN => n10374);
   OUT2_reg_18_inst : DFF_X1 port map( D => n10486, CK => n907, Q => OUT2(18), 
                           QN => n10373);
   OUT2_reg_17_inst : DFF_X1 port map( D => n10489, CK => n903, Q => OUT2(17), 
                           QN => n10372);
   OUT2_reg_16_inst : DFF_X1 port map( D => n10492, CK => n960, Q => OUT2(16), 
                           QN => n10371);
   OUT2_reg_15_inst : DFF_X1 port map( D => n10495, CK => n899, Q => OUT2(15), 
                           QN => n10370);
   OUT2_reg_14_inst : DFF_X1 port map( D => n10498, CK => n876, Q => OUT2(14), 
                           QN => n10369);
   OUT2_reg_13_inst : DFF_X1 port map( D => n10501, CK => n873, Q => OUT2(13), 
                           QN => n10368);
   OUT2_reg_12_inst : DFF_X1 port map( D => n10504, CK => n945, Q => OUT2(12), 
                           QN => n10367);
   OUT2_reg_11_inst : DFF_X1 port map( D => n10507, CK => n880, Q => OUT2(11), 
                           QN => n10366);
   OUT2_reg_10_inst : DFF_X1 port map( D => n10510, CK => n869, Q => OUT2(10), 
                           QN => n10365);
   OUT2_reg_9_inst : DFF_X1 port map( D => n10513, CK => n949, Q => OUT2(9), QN
                           => n10364);
   OUT2_reg_8_inst : DFF_X1 port map( D => n10516, CK => n884, Q => OUT2(8), QN
                           => n10363);
   OUT2_reg_7_inst : DFF_X1 port map( D => n10519, CK => n865, Q => OUT2(7), QN
                           => n10362);
   OUT2_reg_6_inst : DFF_X1 port map( D => n10522, CK => n861, Q => OUT2(6), QN
                           => n10361);
   OUT2_reg_5_inst : DFF_X1 port map( D => n10525, CK => n888, Q => OUT2(5), QN
                           => n10360);
   OUT2_reg_4_inst : DFF_X1 port map( D => n10528, CK => n964, Q => OUT2(4), QN
                           => n10359);
   OUT2_reg_3_inst : DFF_X1 port map( D => n10531, CK => n857, Q => OUT2(3), QN
                           => n10358);
   OUT2_reg_2_inst : DFF_X1 port map( D => n10534, CK => n853, Q => OUT2(2), QN
                           => n10357);
   OUT2_reg_1_inst : DFF_X1 port map( D => n10537, CK => n850, Q => OUT2(1), QN
                           => n10356);
   OUT2_reg_0_inst : DFF_X1 port map( D => n10540, CK => n968, Q => OUT2(0), QN
                           => n10355);
   OUT1_reg_31_inst : DFF_X1 port map( D => n10446, CK => n953, Q => OUT1(31), 
                           QN => n10354);
   OUT1_reg_30_inst : DFF_X1 port map( D => n10449, CK => n895, Q => OUT1(30), 
                           QN => n10353);
   OUT1_reg_29_inst : DFF_X1 port map( D => n10452, CK => n892, Q => OUT1(29), 
                           QN => n10352);
   OUT1_reg_28_inst : DFF_X1 port map( D => n10455, CK => n956, Q => OUT1(28), 
                           QN => n10351);
   OUT1_reg_27_inst : DFF_X1 port map( D => n10458, CK => n937, Q => OUT1(27), 
                           QN => n10350);
   OUT1_reg_26_inst : DFF_X1 port map( D => n10461, CK => n934, Q => OUT1(26), 
                           QN => n10349);
   OUT1_reg_25_inst : DFF_X1 port map( D => n10464, CK => n930, Q => OUT1(25), 
                           QN => n10348);
   OUT1_reg_24_inst : DFF_X1 port map( D => n10467, CK => n941, Q => OUT1(24), 
                           QN => n10347);
   OUT1_reg_23_inst : DFF_X1 port map( D => n10470, CK => n926, Q => OUT1(23), 
                           QN => n10346);
   OUT1_reg_22_inst : DFF_X1 port map( D => n10473, CK => n922, Q => OUT1(22), 
                           QN => n10345);
   OUT1_reg_21_inst : DFF_X1 port map( D => n10476, CK => n918, Q => OUT1(21), 
                           QN => n10344);
   OUT1_reg_20_inst : DFF_X1 port map( D => n10479, CK => n914, Q => OUT1(20), 
                           QN => n10343);
   OUT1_reg_19_inst : DFF_X1 port map( D => n10482, CK => n911, Q => OUT1(19), 
                           QN => n10342);
   OUT1_reg_18_inst : DFF_X1 port map( D => n10485, CK => n907, Q => OUT1(18), 
                           QN => n10341);
   OUT1_reg_17_inst : DFF_X1 port map( D => n10488, CK => n903, Q => OUT1(17), 
                           QN => n10340);
   OUT1_reg_16_inst : DFF_X1 port map( D => n10491, CK => n960, Q => OUT1(16), 
                           QN => n10339);
   OUT1_reg_15_inst : DFF_X1 port map( D => n10494, CK => n899, Q => OUT1(15), 
                           QN => n10338);
   OUT1_reg_14_inst : DFF_X1 port map( D => n10497, CK => n876, Q => OUT1(14), 
                           QN => n10337);
   OUT1_reg_13_inst : DFF_X1 port map( D => n10500, CK => n872, Q => OUT1(13), 
                           QN => n10336);
   OUT1_reg_12_inst : DFF_X1 port map( D => n10503, CK => n945, Q => OUT1(12), 
                           QN => n10335);
   OUT1_reg_11_inst : DFF_X1 port map( D => n10506, CK => n880, Q => OUT1(11), 
                           QN => n10334);
   OUT1_reg_10_inst : DFF_X1 port map( D => n10509, CK => n869, Q => OUT1(10), 
                           QN => n10333);
   OUT1_reg_9_inst : DFF_X1 port map( D => n10512, CK => n949, Q => OUT1(9), QN
                           => n10332);
   OUT1_reg_8_inst : DFF_X1 port map( D => n10515, CK => n884, Q => OUT1(8), QN
                           => n10331);
   OUT1_reg_7_inst : DFF_X1 port map( D => n10518, CK => n865, Q => OUT1(7), QN
                           => n10330);
   OUT1_reg_6_inst : DFF_X1 port map( D => n10521, CK => n861, Q => OUT1(6), QN
                           => n10329);
   OUT1_reg_5_inst : DFF_X1 port map( D => n10524, CK => n888, Q => OUT1(5), QN
                           => n10328);
   OUT1_reg_4_inst : DFF_X1 port map( D => n10527, CK => n964, Q => OUT1(4), QN
                           => n10327);
   OUT1_reg_3_inst : DFF_X1 port map( D => n10530, CK => n857, Q => OUT1(3), QN
                           => n10326);
   OUT1_reg_2_inst : DFF_X1 port map( D => n10533, CK => n853, Q => OUT1(2), QN
                           => n10325);
   OUT1_reg_1_inst : DFF_X1 port map( D => n10536, CK => n850, Q => OUT1(1), QN
                           => n10324);
   OUT1_reg_0_inst : DFF_X1 port map( D => n10539, CK => n972, Q => OUT1(0), QN
                           => n10323);
   REGISTERS_reg_38_30_inst : DFF_X1 port map( D => n13090, CK => n899, Q => 
                           REGISTERS_38_30_port, QN => n11727);
   REGISTERS_reg_39_30_inst : DFF_X1 port map( D => n13122, CK => n899, Q => 
                           REGISTERS_39_30_port, QN => n11759);
   REGISTERS_reg_37_30_inst : DFF_X1 port map( D => n13058, CK => n899, Q => 
                           REGISTERS_37_30_port, QN => n11695);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n11874, CK => n899, Q => 
                           REGISTERS_0_30_port, QN => n10451);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n11906, CK => n899, Q => 
                           REGISTERS_1_30_port, QN => n10543);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n11938, CK => n899, Q => 
                           REGISTERS_2_30_port, QN => n10575);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n11970, CK => n898, Q => 
                           REGISTERS_3_30_port, QN => n10607);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n12002, CK => n898, Q => 
                           REGISTERS_4_30_port, QN => n10639);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n12034, CK => n898, Q => 
                           REGISTERS_5_30_port, QN => n10671);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n12066, CK => n898, Q => 
                           REGISTERS_6_30_port, QN => n10703);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n12098, CK => n898, Q => 
                           REGISTERS_7_30_port, QN => n10735);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n12130, CK => n898, Q => 
                           REGISTERS_8_30_port, QN => n10767);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n12162, CK => n898, Q => 
                           REGISTERS_9_30_port, QN => n10799);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n12194, CK => n898, Q => 
                           REGISTERS_10_30_port, QN => n10831);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n12226_port, CK => n898, Q 
                           => REGISTERS_11_30_port, QN => n10863);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n12258_port, CK => n898, Q 
                           => REGISTERS_12_30_port, QN => n10895);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n12290_port, CK => n898, Q 
                           => REGISTERS_13_30_port, QN => n10927);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n12322, CK => n897, Q => 
                           REGISTERS_14_30_port, QN => n10959);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n12354, CK => n897, Q => 
                           REGISTERS_15_30_port, QN => n10991);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n12386, CK => n897, Q => 
                           REGISTERS_16_30_port, QN => n11023);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n12418, CK => n897, Q => 
                           REGISTERS_17_30_port, QN => n11055);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n12450, CK => n897, Q => 
                           REGISTERS_18_30_port, QN => n11087);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n12482, CK => n897, Q => 
                           REGISTERS_19_30_port, QN => n11119);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n12514, CK => n897, Q => 
                           REGISTERS_20_30_port, QN => n11151);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n12546, CK => n897, Q => 
                           REGISTERS_21_30_port, QN => n11183);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n12578, CK => n897, Q => 
                           REGISTERS_22_30_port, QN => n11215);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n12610, CK => n897, Q => 
                           REGISTERS_23_30_port, QN => n11247);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n12642, CK => n897, Q => 
                           REGISTERS_24_30_port, QN => n11279);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n12674, CK => n896, Q => 
                           REGISTERS_25_30_port, QN => n11311);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n12706, CK => n896, Q => 
                           REGISTERS_26_30_port, QN => n11343);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n12738, CK => n896, Q => 
                           REGISTERS_27_30_port, QN => n11375);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n12770, CK => n896, Q => 
                           REGISTERS_28_30_port, QN => n11407);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n12802, CK => n896, Q => 
                           REGISTERS_29_30_port, QN => n11439);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n12834, CK => n896, Q => 
                           REGISTERS_30_30_port, QN => n11471);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n12866, CK => n896, Q => 
                           REGISTERS_31_30_port, QN => n11503);
   REGISTERS_reg_32_30_inst : DFF_X1 port map( D => n12898, CK => n896, Q => 
                           REGISTERS_32_30_port, QN => n11535);
   REGISTERS_reg_33_30_inst : DFF_X1 port map( D => n12930, CK => n896, Q => 
                           REGISTERS_33_30_port, QN => n11567);
   REGISTERS_reg_34_30_inst : DFF_X1 port map( D => n12962, CK => n896, Q => 
                           REGISTERS_34_30_port, QN => n11599);
   REGISTERS_reg_35_30_inst : DFF_X1 port map( D => n12994, CK => n896, Q => 
                           REGISTERS_35_30_port, QN => n11631);
   REGISTERS_reg_36_30_inst : DFF_X1 port map( D => n13026, CK => n899, Q => 
                           REGISTERS_36_30_port, QN => n11663);
   REGISTERS_reg_38_29_inst : DFF_X1 port map( D => n13091, CK => n895, Q => 
                           REGISTERS_38_29_port, QN => n11728);
   REGISTERS_reg_39_29_inst : DFF_X1 port map( D => n13123, CK => n895, Q => 
                           REGISTERS_39_29_port, QN => n11760);
   REGISTERS_reg_37_29_inst : DFF_X1 port map( D => n13059, CK => n895, Q => 
                           REGISTERS_37_29_port, QN => n11696);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n11875, CK => n895, Q => 
                           REGISTERS_0_29_port, QN => n10454);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n11907, CK => n895, Q => 
                           REGISTERS_1_29_port, QN => n10544);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n11939, CK => n895, Q => 
                           REGISTERS_2_29_port, QN => n10576);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n11971, CK => n895, Q => 
                           REGISTERS_3_29_port, QN => n10608);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n12003, CK => n895, Q => 
                           REGISTERS_4_29_port, QN => n10640);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n12035, CK => n894, Q => 
                           REGISTERS_5_29_port, QN => n10672);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n12067, CK => n894, Q => 
                           REGISTERS_6_29_port, QN => n10704);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n12099, CK => n894, Q => 
                           REGISTERS_7_29_port, QN => n10736);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n12131, CK => n894, Q => 
                           REGISTERS_8_29_port, QN => n10768);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n12163, CK => n894, Q => 
                           REGISTERS_9_29_port, QN => n10800);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n12195, CK => n894, Q => 
                           REGISTERS_10_29_port, QN => n10832);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n12227_port, CK => n894, Q 
                           => REGISTERS_11_29_port, QN => n10864);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n12259_port, CK => n894, Q 
                           => REGISTERS_12_29_port, QN => n10896);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n12291_port, CK => n894, Q 
                           => REGISTERS_13_29_port, QN => n10928);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n12323, CK => n894, Q => 
                           REGISTERS_14_29_port, QN => n10960);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n12355, CK => n894, Q => 
                           REGISTERS_15_29_port, QN => n10992);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n12387, CK => n893, Q => 
                           REGISTERS_16_29_port, QN => n11024);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n12419, CK => n893, Q => 
                           REGISTERS_17_29_port, QN => n11056);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n12451, CK => n893, Q => 
                           REGISTERS_18_29_port, QN => n11088);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n12483, CK => n893, Q => 
                           REGISTERS_19_29_port, QN => n11120);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n12515, CK => n893, Q => 
                           REGISTERS_20_29_port, QN => n11152);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n12547, CK => n893, Q => 
                           REGISTERS_21_29_port, QN => n11184);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n12579, CK => n893, Q => 
                           REGISTERS_22_29_port, QN => n11216);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n12611, CK => n893, Q => 
                           REGISTERS_23_29_port, QN => n11248);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n12643, CK => n893, Q => 
                           REGISTERS_24_29_port, QN => n11280);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n12675, CK => n893, Q => 
                           REGISTERS_25_29_port, QN => n11312);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n12707, CK => n893, Q => 
                           REGISTERS_26_29_port, QN => n11344);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n12739, CK => n892, Q => 
                           REGISTERS_27_29_port, QN => n11376);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n12771, CK => n892, Q => 
                           REGISTERS_28_29_port, QN => n11408);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n12803, CK => n892, Q => 
                           REGISTERS_29_29_port, QN => n11440);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n12835, CK => n892, Q => 
                           REGISTERS_30_29_port, QN => n11472);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n12867, CK => n892, Q => 
                           REGISTERS_31_29_port, QN => n11504);
   REGISTERS_reg_32_29_inst : DFF_X1 port map( D => n12899, CK => n892, Q => 
                           REGISTERS_32_29_port, QN => n11536);
   REGISTERS_reg_33_29_inst : DFF_X1 port map( D => n12931, CK => n892, Q => 
                           REGISTERS_33_29_port, QN => n11568);
   REGISTERS_reg_34_29_inst : DFF_X1 port map( D => n12963, CK => n892, Q => 
                           REGISTERS_34_29_port, QN => n11600);
   REGISTERS_reg_35_29_inst : DFF_X1 port map( D => n12995, CK => n892, Q => 
                           REGISTERS_35_29_port, QN => n11632);
   REGISTERS_reg_36_29_inst : DFF_X1 port map( D => n13027, CK => n895, Q => 
                           REGISTERS_36_29_port, QN => n11664);
   REGISTERS_reg_38_28_inst : DFF_X1 port map( D => n13092, CK => n960, Q => 
                           REGISTERS_38_28_port, QN => n11729);
   REGISTERS_reg_39_28_inst : DFF_X1 port map( D => n13124, CK => n960, Q => 
                           REGISTERS_39_28_port, QN => n11761);
   REGISTERS_reg_37_28_inst : DFF_X1 port map( D => n13060, CK => n960, Q => 
                           REGISTERS_37_28_port, QN => n11697);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n11876, CK => n960, Q => 
                           REGISTERS_0_28_port, QN => n10457);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n11908, CK => n960, Q => 
                           REGISTERS_1_28_port, QN => n10545);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n11940, CK => n960, Q => 
                           REGISTERS_2_28_port, QN => n10577);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n11972, CK => n960, Q => 
                           REGISTERS_3_28_port, QN => n10609);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n12004, CK => n959, Q => 
                           REGISTERS_4_28_port, QN => n10641);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n12036, CK => n959, Q => 
                           REGISTERS_5_28_port, QN => n10673);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n12068, CK => n959, Q => 
                           REGISTERS_6_28_port, QN => n10705);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n12100, CK => n959, Q => 
                           REGISTERS_7_28_port, QN => n10737);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n12132, CK => n959, Q => 
                           REGISTERS_8_28_port, QN => n10769);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n12164, CK => n959, Q => 
                           REGISTERS_9_28_port, QN => n10801);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n12196, CK => n959, Q => 
                           REGISTERS_10_28_port, QN => n10833);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n12228_port, CK => n959, Q 
                           => REGISTERS_11_28_port, QN => n10865);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n12260_port, CK => n959, Q 
                           => REGISTERS_12_28_port, QN => n10897);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n12292_port, CK => n959, Q 
                           => REGISTERS_13_28_port, QN => n10929);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n12324, CK => n959, Q => 
                           REGISTERS_14_28_port, QN => n10961);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n12356, CK => n958, Q => 
                           REGISTERS_15_28_port, QN => n10993);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n12388, CK => n958, Q => 
                           REGISTERS_16_28_port, QN => n11025);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n12420, CK => n958, Q => 
                           REGISTERS_17_28_port, QN => n11057);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n12452, CK => n958, Q => 
                           REGISTERS_18_28_port, QN => n11089);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n12484, CK => n958, Q => 
                           REGISTERS_19_28_port, QN => n11121);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n12516, CK => n958, Q => 
                           REGISTERS_20_28_port, QN => n11153);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n12548, CK => n958, Q => 
                           REGISTERS_21_28_port, QN => n11185);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n12580, CK => n958, Q => 
                           REGISTERS_22_28_port, QN => n11217);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n12612, CK => n958, Q => 
                           REGISTERS_23_28_port, QN => n11249);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n12644, CK => n958, Q => 
                           REGISTERS_24_28_port, QN => n11281);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n12676, CK => n958, Q => 
                           REGISTERS_25_28_port, QN => n11313);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n12708, CK => n957, Q => 
                           REGISTERS_26_28_port, QN => n11345);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n12740, CK => n957, Q => 
                           REGISTERS_27_28_port, QN => n11377);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n12772, CK => n957, Q => 
                           REGISTERS_28_28_port, QN => n11409);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n12804, CK => n957, Q => 
                           REGISTERS_29_28_port, QN => n11441);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n12836, CK => n957, Q => 
                           REGISTERS_30_28_port, QN => n11473);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n12868, CK => n957, Q => 
                           REGISTERS_31_28_port, QN => n11505);
   REGISTERS_reg_32_28_inst : DFF_X1 port map( D => n12900, CK => n957, Q => 
                           REGISTERS_32_28_port, QN => n11537);
   REGISTERS_reg_33_28_inst : DFF_X1 port map( D => n12932, CK => n957, Q => 
                           REGISTERS_33_28_port, QN => n11569);
   REGISTERS_reg_34_28_inst : DFF_X1 port map( D => n12964, CK => n957, Q => 
                           REGISTERS_34_28_port, QN => n11601);
   REGISTERS_reg_35_28_inst : DFF_X1 port map( D => n12996, CK => n957, Q => 
                           REGISTERS_35_28_port, QN => n11633);
   REGISTERS_reg_36_28_inst : DFF_X1 port map( D => n13028, CK => n960, Q => 
                           REGISTERS_36_28_port, QN => n11665);
   REGISTERS_reg_38_27_inst : DFF_X1 port map( D => n13093, CK => n941, Q => 
                           REGISTERS_38_27_port, QN => n11730);
   REGISTERS_reg_39_27_inst : DFF_X1 port map( D => n13125, CK => n941, Q => 
                           REGISTERS_39_27_port, QN => n11762);
   REGISTERS_reg_37_27_inst : DFF_X1 port map( D => n13061, CK => n941, Q => 
                           REGISTERS_37_27_port, QN => n11698);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n11877, CK => n941, Q => 
                           REGISTERS_0_27_port, QN => n10460);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n11909, CK => n941, Q => 
                           REGISTERS_1_27_port, QN => n10546);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n11941, CK => n941, Q => 
                           REGISTERS_2_27_port, QN => n10578);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n11973, CK => n940, Q => 
                           REGISTERS_3_27_port, QN => n10610);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n12005, CK => n940, Q => 
                           REGISTERS_4_27_port, QN => n10642);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n12037, CK => n940, Q => 
                           REGISTERS_5_27_port, QN => n10674);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n12069, CK => n940, Q => 
                           REGISTERS_6_27_port, QN => n10706);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n12101, CK => n940, Q => 
                           REGISTERS_7_27_port, QN => n10738);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n12133, CK => n940, Q => 
                           REGISTERS_8_27_port, QN => n10770);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n12165, CK => n940, Q => 
                           REGISTERS_9_27_port, QN => n10802);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n12197, CK => n940, Q => 
                           REGISTERS_10_27_port, QN => n10834);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n12229_port, CK => n940, Q 
                           => REGISTERS_11_27_port, QN => n10866);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n12261_port, CK => n940, Q 
                           => REGISTERS_12_27_port, QN => n10898);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n12293_port, CK => n940, Q 
                           => REGISTERS_13_27_port, QN => n10930);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n12325, CK => n939, Q => 
                           REGISTERS_14_27_port, QN => n10962);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n12357, CK => n939, Q => 
                           REGISTERS_15_27_port, QN => n10994);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n12389, CK => n939, Q => 
                           REGISTERS_16_27_port, QN => n11026);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n12421, CK => n939, Q => 
                           REGISTERS_17_27_port, QN => n11058);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n12453, CK => n939, Q => 
                           REGISTERS_18_27_port, QN => n11090);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n12485, CK => n939, Q => 
                           REGISTERS_19_27_port, QN => n11122);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n12517, CK => n939, Q => 
                           REGISTERS_20_27_port, QN => n11154);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n12549, CK => n939, Q => 
                           REGISTERS_21_27_port, QN => n11186);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n12581, CK => n939, Q => 
                           REGISTERS_22_27_port, QN => n11218);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n12613, CK => n939, Q => 
                           REGISTERS_23_27_port, QN => n11250);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n12645, CK => n939, Q => 
                           REGISTERS_24_27_port, QN => n11282);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n12677, CK => n938, Q => 
                           REGISTERS_25_27_port, QN => n11314);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n12709, CK => n938, Q => 
                           REGISTERS_26_27_port, QN => n11346);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n12741, CK => n938, Q => 
                           REGISTERS_27_27_port, QN => n11378);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n12773, CK => n938, Q => 
                           REGISTERS_28_27_port, QN => n11410);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n12805, CK => n938, Q => 
                           REGISTERS_29_27_port, QN => n11442);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n12837, CK => n938, Q => 
                           REGISTERS_30_27_port, QN => n11474);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n12869, CK => n938, Q => 
                           REGISTERS_31_27_port, QN => n11506);
   REGISTERS_reg_32_27_inst : DFF_X1 port map( D => n12901, CK => n938, Q => 
                           REGISTERS_32_27_port, QN => n11538);
   REGISTERS_reg_33_27_inst : DFF_X1 port map( D => n12933, CK => n938, Q => 
                           REGISTERS_33_27_port, QN => n11570);
   REGISTERS_reg_34_27_inst : DFF_X1 port map( D => n12965, CK => n938, Q => 
                           REGISTERS_34_27_port, QN => n11602);
   REGISTERS_reg_35_27_inst : DFF_X1 port map( D => n12997, CK => n938, Q => 
                           REGISTERS_35_27_port, QN => n11634);
   REGISTERS_reg_36_27_inst : DFF_X1 port map( D => n13029, CK => n941, Q => 
                           REGISTERS_36_27_port, QN => n11666);
   REGISTERS_reg_38_26_inst : DFF_X1 port map( D => n13094, CK => n937, Q => 
                           REGISTERS_38_26_port, QN => n11731);
   REGISTERS_reg_39_26_inst : DFF_X1 port map( D => n13126, CK => n937, Q => 
                           REGISTERS_39_26_port, QN => n11763);
   REGISTERS_reg_37_26_inst : DFF_X1 port map( D => n13062, CK => n937, Q => 
                           REGISTERS_37_26_port, QN => n11699);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n11878, CK => n937, Q => 
                           REGISTERS_0_26_port, QN => n10463);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n11910, CK => n937, Q => 
                           REGISTERS_1_26_port, QN => n10547);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n11942, CK => n937, Q => 
                           REGISTERS_2_26_port, QN => n10579);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n11974, CK => n937, Q => 
                           REGISTERS_3_26_port, QN => n10611);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n12006, CK => n937, Q => 
                           REGISTERS_4_26_port, QN => n10643);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n12038, CK => n936, Q => 
                           REGISTERS_5_26_port, QN => n10675);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n12070, CK => n936, Q => 
                           REGISTERS_6_26_port, QN => n10707);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n12102, CK => n936, Q => 
                           REGISTERS_7_26_port, QN => n10739);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n12134, CK => n936, Q => 
                           REGISTERS_8_26_port, QN => n10771);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n12166, CK => n936, Q => 
                           REGISTERS_9_26_port, QN => n10803);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n12198, CK => n936, Q => 
                           REGISTERS_10_26_port, QN => n10835);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n12230_port, CK => n936, Q 
                           => REGISTERS_11_26_port, QN => n10867);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n12262_port, CK => n936, Q 
                           => REGISTERS_12_26_port, QN => n10899);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n12294_port, CK => n936, Q 
                           => REGISTERS_13_26_port, QN => n10931);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n12326, CK => n936, Q => 
                           REGISTERS_14_26_port, QN => n10963);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n12358, CK => n936, Q => 
                           REGISTERS_15_26_port, QN => n10995);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n12390, CK => n935, Q => 
                           REGISTERS_16_26_port, QN => n11027);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n12422, CK => n935, Q => 
                           REGISTERS_17_26_port, QN => n11059);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n12454, CK => n935, Q => 
                           REGISTERS_18_26_port, QN => n11091);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n12486, CK => n935, Q => 
                           REGISTERS_19_26_port, QN => n11123);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n12518, CK => n935, Q => 
                           REGISTERS_20_26_port, QN => n11155);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n12550, CK => n935, Q => 
                           REGISTERS_21_26_port, QN => n11187);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n12582, CK => n935, Q => 
                           REGISTERS_22_26_port, QN => n11219);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n12614, CK => n935, Q => 
                           REGISTERS_23_26_port, QN => n11251);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n12646, CK => n935, Q => 
                           REGISTERS_24_26_port, QN => n11283);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n12678, CK => n935, Q => 
                           REGISTERS_25_26_port, QN => n11315);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n12710, CK => n935, Q => 
                           REGISTERS_26_26_port, QN => n11347);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n12742, CK => n934, Q => 
                           REGISTERS_27_26_port, QN => n11379);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n12774, CK => n934, Q => 
                           REGISTERS_28_26_port, QN => n11411);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n12806, CK => n934, Q => 
                           REGISTERS_29_26_port, QN => n11443);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n12838, CK => n934, Q => 
                           REGISTERS_30_26_port, QN => n11475);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n12870, CK => n934, Q => 
                           REGISTERS_31_26_port, QN => n11507);
   REGISTERS_reg_32_26_inst : DFF_X1 port map( D => n12902, CK => n934, Q => 
                           REGISTERS_32_26_port, QN => n11539);
   REGISTERS_reg_33_26_inst : DFF_X1 port map( D => n12934, CK => n934, Q => 
                           REGISTERS_33_26_port, QN => n11571);
   REGISTERS_reg_34_26_inst : DFF_X1 port map( D => n12966, CK => n934, Q => 
                           REGISTERS_34_26_port, QN => n11603);
   REGISTERS_reg_35_26_inst : DFF_X1 port map( D => n12998, CK => n934, Q => 
                           REGISTERS_35_26_port, QN => n11635);
   REGISTERS_reg_36_26_inst : DFF_X1 port map( D => n13030, CK => n937, Q => 
                           REGISTERS_36_26_port, QN => n11667);
   REGISTERS_reg_38_25_inst : DFF_X1 port map( D => n13095, CK => n933, Q => 
                           REGISTERS_38_25_port, QN => n11732);
   REGISTERS_reg_39_25_inst : DFF_X1 port map( D => n13127, CK => n933, Q => 
                           REGISTERS_39_25_port, QN => n11764);
   REGISTERS_reg_37_25_inst : DFF_X1 port map( D => n13063, CK => n933, Q => 
                           REGISTERS_37_25_port, QN => n11700);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n11879, CK => n933, Q => 
                           REGISTERS_0_25_port, QN => n10466);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n11911, CK => n933, Q => 
                           REGISTERS_1_25_port, QN => n10548);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n11943, CK => n933, Q => 
                           REGISTERS_2_25_port, QN => n10580);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n11975, CK => n933, Q => 
                           REGISTERS_3_25_port, QN => n10612);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n12007, CK => n933, Q => 
                           REGISTERS_4_25_port, QN => n10644);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n12039, CK => n933, Q => 
                           REGISTERS_5_25_port, QN => n10676);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n12071, CK => n933, Q => 
                           REGISTERS_6_25_port, QN => n10708);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n12103, CK => n932, Q => 
                           REGISTERS_7_25_port, QN => n10740);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n12135, CK => n932, Q => 
                           REGISTERS_8_25_port, QN => n10772);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n12167, CK => n932, Q => 
                           REGISTERS_9_25_port, QN => n10804);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n12199, CK => n932, Q => 
                           REGISTERS_10_25_port, QN => n10836);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n12231_port, CK => n932, Q 
                           => REGISTERS_11_25_port, QN => n10868);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n12263_port, CK => n932, Q 
                           => REGISTERS_12_25_port, QN => n10900);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n12295_port, CK => n932, Q 
                           => REGISTERS_13_25_port, QN => n10932);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n12327, CK => n932, Q => 
                           REGISTERS_14_25_port, QN => n10964);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n12359, CK => n932, Q => 
                           REGISTERS_15_25_port, QN => n10996);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n12391, CK => n932, Q => 
                           REGISTERS_16_25_port, QN => n11028);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n12423, CK => n932, Q => 
                           REGISTERS_17_25_port, QN => n11060);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n12455, CK => n931, Q => 
                           REGISTERS_18_25_port, QN => n11092);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n12487, CK => n931, Q => 
                           REGISTERS_19_25_port, QN => n11124);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n12519, CK => n931, Q => 
                           REGISTERS_20_25_port, QN => n11156);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n12551, CK => n931, Q => 
                           REGISTERS_21_25_port, QN => n11188);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n12583, CK => n931, Q => 
                           REGISTERS_22_25_port, QN => n11220);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n12615, CK => n931, Q => 
                           REGISTERS_23_25_port, QN => n11252);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n12647, CK => n931, Q => 
                           REGISTERS_24_25_port, QN => n11284);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n12679, CK => n931, Q => 
                           REGISTERS_25_25_port, QN => n11316);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n12711, CK => n931, Q => 
                           REGISTERS_26_25_port, QN => n11348);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n12743, CK => n931, Q => 
                           REGISTERS_27_25_port, QN => n11380);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n12775, CK => n931, Q => 
                           REGISTERS_28_25_port, QN => n11412);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n12807, CK => n930, Q => 
                           REGISTERS_29_25_port, QN => n11444);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n12839, CK => n930, Q => 
                           REGISTERS_30_25_port, QN => n11476);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n12871, CK => n930, Q => 
                           REGISTERS_31_25_port, QN => n11508);
   REGISTERS_reg_32_25_inst : DFF_X1 port map( D => n12903, CK => n930, Q => 
                           REGISTERS_32_25_port, QN => n11540);
   REGISTERS_reg_33_25_inst : DFF_X1 port map( D => n12935, CK => n930, Q => 
                           REGISTERS_33_25_port, QN => n11572);
   REGISTERS_reg_34_25_inst : DFF_X1 port map( D => n12967, CK => n930, Q => 
                           REGISTERS_34_25_port, QN => n11604);
   REGISTERS_reg_35_25_inst : DFF_X1 port map( D => n12999, CK => n930, Q => 
                           REGISTERS_35_25_port, QN => n11636);
   REGISTERS_reg_36_25_inst : DFF_X1 port map( D => n13031, CK => n933, Q => 
                           REGISTERS_36_25_port, QN => n11668);
   REGISTERS_reg_38_24_inst : DFF_X1 port map( D => n13096, CK => n945, Q => 
                           REGISTERS_38_24_port, QN => n11733);
   REGISTERS_reg_39_24_inst : DFF_X1 port map( D => n13128, CK => n945, Q => 
                           REGISTERS_39_24_port, QN => n11765);
   REGISTERS_reg_37_24_inst : DFF_X1 port map( D => n13064, CK => n945, Q => 
                           REGISTERS_37_24_port, QN => n11701);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n11880, CK => n945, Q => 
                           REGISTERS_0_24_port, QN => n10469);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n11912, CK => n944, Q => 
                           REGISTERS_1_24_port, QN => n10549);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n11944, CK => n944, Q => 
                           REGISTERS_2_24_port, QN => n10581);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n11976, CK => n944, Q => 
                           REGISTERS_3_24_port, QN => n10613);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n12008, CK => n944, Q => 
                           REGISTERS_4_24_port, QN => n10645);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n12040, CK => n944, Q => 
                           REGISTERS_5_24_port, QN => n10677);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n12072, CK => n944, Q => 
                           REGISTERS_6_24_port, QN => n10709);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n12104, CK => n944, Q => 
                           REGISTERS_7_24_port, QN => n10741);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n12136, CK => n944, Q => 
                           REGISTERS_8_24_port, QN => n10773);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n12168, CK => n944, Q => 
                           REGISTERS_9_24_port, QN => n10805);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n12200, CK => n944, Q => 
                           REGISTERS_10_24_port, QN => n10837);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n12232_port, CK => n944, Q 
                           => REGISTERS_11_24_port, QN => n10869);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n12264_port, CK => n943, Q 
                           => REGISTERS_12_24_port, QN => n10901);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n12296_port, CK => n943, Q 
                           => REGISTERS_13_24_port, QN => n10933);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n12328, CK => n943, Q => 
                           REGISTERS_14_24_port, QN => n10965);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n12360, CK => n943, Q => 
                           REGISTERS_15_24_port, QN => n10997);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n12392, CK => n943, Q => 
                           REGISTERS_16_24_port, QN => n11029);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n12424, CK => n943, Q => 
                           REGISTERS_17_24_port, QN => n11061);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n12456, CK => n943, Q => 
                           REGISTERS_18_24_port, QN => n11093);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n12488, CK => n943, Q => 
                           REGISTERS_19_24_port, QN => n11125);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n12520, CK => n943, Q => 
                           REGISTERS_20_24_port, QN => n11157);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n12552, CK => n943, Q => 
                           REGISTERS_21_24_port, QN => n11189);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n12584, CK => n943, Q => 
                           REGISTERS_22_24_port, QN => n11221);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n12616, CK => n942, Q => 
                           REGISTERS_23_24_port, QN => n11253);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n12648, CK => n942, Q => 
                           REGISTERS_24_24_port, QN => n11285);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n12680, CK => n942, Q => 
                           REGISTERS_25_24_port, QN => n11317);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n12712, CK => n942, Q => 
                           REGISTERS_26_24_port, QN => n11349);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n12744, CK => n942, Q => 
                           REGISTERS_27_24_port, QN => n11381);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n12776, CK => n942, Q => 
                           REGISTERS_28_24_port, QN => n11413);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n12808, CK => n942, Q => 
                           REGISTERS_29_24_port, QN => n11445);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n12840, CK => n942, Q => 
                           REGISTERS_30_24_port, QN => n11477);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n12872, CK => n942, Q => 
                           REGISTERS_31_24_port, QN => n11509);
   REGISTERS_reg_32_24_inst : DFF_X1 port map( D => n12904, CK => n942, Q => 
                           REGISTERS_32_24_port, QN => n11541);
   REGISTERS_reg_33_24_inst : DFF_X1 port map( D => n12936, CK => n942, Q => 
                           REGISTERS_33_24_port, QN => n11573);
   REGISTERS_reg_34_24_inst : DFF_X1 port map( D => n12968, CK => n941, Q => 
                           REGISTERS_34_24_port, QN => n11605);
   REGISTERS_reg_35_24_inst : DFF_X1 port map( D => n13000, CK => n941, Q => 
                           REGISTERS_35_24_port, QN => n11637);
   REGISTERS_reg_36_24_inst : DFF_X1 port map( D => n13032, CK => n945, Q => 
                           REGISTERS_36_24_port, QN => n11669);
   REGISTERS_reg_38_23_inst : DFF_X1 port map( D => n13097, CK => n929, Q => 
                           REGISTERS_38_23_port, QN => n11734);
   REGISTERS_reg_39_23_inst : DFF_X1 port map( D => n13129, CK => n930, Q => 
                           REGISTERS_39_23_port, QN => n11766);
   REGISTERS_reg_37_23_inst : DFF_X1 port map( D => n13065, CK => n929, Q => 
                           REGISTERS_37_23_port, QN => n11702);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n11881, CK => n929, Q => 
                           REGISTERS_0_23_port, QN => n10472);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n11913, CK => n929, Q => 
                           REGISTERS_1_23_port, QN => n10550);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n11945, CK => n929, Q => 
                           REGISTERS_2_23_port, QN => n10582);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n11977, CK => n929, Q => 
                           REGISTERS_3_23_port, QN => n10614);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n12009, CK => n929, Q => 
                           REGISTERS_4_23_port, QN => n10646);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n12041, CK => n929, Q => 
                           REGISTERS_5_23_port, QN => n10678);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n12073, CK => n929, Q => 
                           REGISTERS_6_23_port, QN => n10710);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n12105, CK => n929, Q => 
                           REGISTERS_7_23_port, QN => n10742);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n12137, CK => n929, Q => 
                           REGISTERS_8_23_port, QN => n10774);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n12169, CK => n928, Q => 
                           REGISTERS_9_23_port, QN => n10806);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n12201, CK => n928, Q => 
                           REGISTERS_10_23_port, QN => n10838);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n12233_port, CK => n928, Q 
                           => REGISTERS_11_23_port, QN => n10870);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n12265_port, CK => n928, Q 
                           => REGISTERS_12_23_port, QN => n10902);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n12297_port, CK => n928, Q 
                           => REGISTERS_13_23_port, QN => n10934);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n12329, CK => n928, Q => 
                           REGISTERS_14_23_port, QN => n10966);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n12361, CK => n928, Q => 
                           REGISTERS_15_23_port, QN => n10998);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n12393, CK => n928, Q => 
                           REGISTERS_16_23_port, QN => n11030);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n12425, CK => n928, Q => 
                           REGISTERS_17_23_port, QN => n11062);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n12457, CK => n928, Q => 
                           REGISTERS_18_23_port, QN => n11094);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n12489, CK => n928, Q => 
                           REGISTERS_19_23_port, QN => n11126);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n12521, CK => n927, Q => 
                           REGISTERS_20_23_port, QN => n11158);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n12553, CK => n927, Q => 
                           REGISTERS_21_23_port, QN => n11190);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n12585, CK => n927, Q => 
                           REGISTERS_22_23_port, QN => n11222);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n12617, CK => n927, Q => 
                           REGISTERS_23_23_port, QN => n11254);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n12649, CK => n927, Q => 
                           REGISTERS_24_23_port, QN => n11286);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n12681, CK => n927, Q => 
                           REGISTERS_25_23_port, QN => n11318);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n12713, CK => n927, Q => 
                           REGISTERS_26_23_port, QN => n11350);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n12745, CK => n927, Q => 
                           REGISTERS_27_23_port, QN => n11382);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n12777, CK => n927, Q => 
                           REGISTERS_28_23_port, QN => n11414);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n12809, CK => n927, Q => 
                           REGISTERS_29_23_port, QN => n11446);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n12841, CK => n927, Q => 
                           REGISTERS_30_23_port, QN => n11478);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n12873, CK => n926, Q => 
                           REGISTERS_31_23_port, QN => n11510);
   REGISTERS_reg_32_23_inst : DFF_X1 port map( D => n12905, CK => n926, Q => 
                           REGISTERS_32_23_port, QN => n11542);
   REGISTERS_reg_33_23_inst : DFF_X1 port map( D => n12937, CK => n926, Q => 
                           REGISTERS_33_23_port, QN => n11574);
   REGISTERS_reg_34_23_inst : DFF_X1 port map( D => n12969, CK => n926, Q => 
                           REGISTERS_34_23_port, QN => n11606);
   REGISTERS_reg_35_23_inst : DFF_X1 port map( D => n13001, CK => n926, Q => 
                           REGISTERS_35_23_port, QN => n11638);
   REGISTERS_reg_36_23_inst : DFF_X1 port map( D => n13033, CK => n930, Q => 
                           REGISTERS_36_23_port, QN => n11670);
   REGISTERS_reg_38_22_inst : DFF_X1 port map( D => n13098, CK => n926, Q => 
                           REGISTERS_38_22_port, QN => n11735);
   REGISTERS_reg_39_22_inst : DFF_X1 port map( D => n13130, CK => n926, Q => 
                           REGISTERS_39_22_port, QN => n11767);
   REGISTERS_reg_37_22_inst : DFF_X1 port map( D => n13066, CK => n926, Q => 
                           REGISTERS_37_22_port, QN => n11703);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n11882, CK => n925, Q => 
                           REGISTERS_0_22_port, QN => n10475);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n11914, CK => n925, Q => 
                           REGISTERS_1_22_port, QN => n10551);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n11946, CK => n925, Q => 
                           REGISTERS_2_22_port, QN => n10583);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n11978, CK => n925, Q => 
                           REGISTERS_3_22_port, QN => n10615);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n12010, CK => n925, Q => 
                           REGISTERS_4_22_port, QN => n10647);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n12042, CK => n925, Q => 
                           REGISTERS_5_22_port, QN => n10679);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n12074, CK => n925, Q => 
                           REGISTERS_6_22_port, QN => n10711);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n12106, CK => n925, Q => 
                           REGISTERS_7_22_port, QN => n10743);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n12138, CK => n925, Q => 
                           REGISTERS_8_22_port, QN => n10775);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n12170, CK => n925, Q => 
                           REGISTERS_9_22_port, QN => n10807);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n12202, CK => n925, Q => 
                           REGISTERS_10_22_port, QN => n10839);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n12234_port, CK => n924, Q 
                           => REGISTERS_11_22_port, QN => n10871);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n12266_port, CK => n924, Q 
                           => REGISTERS_12_22_port, QN => n10903);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n12298_port, CK => n924, Q 
                           => REGISTERS_13_22_port, QN => n10935);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n12330, CK => n924, Q => 
                           REGISTERS_14_22_port, QN => n10967);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n12362, CK => n924, Q => 
                           REGISTERS_15_22_port, QN => n10999);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n12394, CK => n924, Q => 
                           REGISTERS_16_22_port, QN => n11031);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n12426, CK => n924, Q => 
                           REGISTERS_17_22_port, QN => n11063);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n12458, CK => n924, Q => 
                           REGISTERS_18_22_port, QN => n11095);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n12490, CK => n924, Q => 
                           REGISTERS_19_22_port, QN => n11127);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n12522, CK => n924, Q => 
                           REGISTERS_20_22_port, QN => n11159);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n12554, CK => n924, Q => 
                           REGISTERS_21_22_port, QN => n11191);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n12586, CK => n923, Q => 
                           REGISTERS_22_22_port, QN => n11223);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n12618, CK => n923, Q => 
                           REGISTERS_23_22_port, QN => n11255);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n12650, CK => n923, Q => 
                           REGISTERS_24_22_port, QN => n11287);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n12682, CK => n923, Q => 
                           REGISTERS_25_22_port, QN => n11319);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n12714, CK => n923, Q => 
                           REGISTERS_26_22_port, QN => n11351);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n12746, CK => n923, Q => 
                           REGISTERS_27_22_port, QN => n11383);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n12778, CK => n923, Q => 
                           REGISTERS_28_22_port, QN => n11415);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n12810, CK => n923, Q => 
                           REGISTERS_29_22_port, QN => n11447);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n12842, CK => n923, Q => 
                           REGISTERS_30_22_port, QN => n11479);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n12874, CK => n923, Q => 
                           REGISTERS_31_22_port, QN => n11511);
   REGISTERS_reg_32_22_inst : DFF_X1 port map( D => n12906, CK => n923, Q => 
                           REGISTERS_32_22_port, QN => n11543);
   REGISTERS_reg_33_22_inst : DFF_X1 port map( D => n12938, CK => n922, Q => 
                           REGISTERS_33_22_port, QN => n11575);
   REGISTERS_reg_34_22_inst : DFF_X1 port map( D => n12970, CK => n922, Q => 
                           REGISTERS_34_22_port, QN => n11607);
   REGISTERS_reg_35_22_inst : DFF_X1 port map( D => n13002, CK => n922, Q => 
                           REGISTERS_35_22_port, QN => n11639);
   REGISTERS_reg_36_22_inst : DFF_X1 port map( D => n13034, CK => n926, Q => 
                           REGISTERS_36_22_port, QN => n11671);
   REGISTERS_reg_38_21_inst : DFF_X1 port map( D => n13099, CK => n922, Q => 
                           REGISTERS_38_21_port, QN => n11736);
   REGISTERS_reg_39_21_inst : DFF_X1 port map( D => n13131, CK => n922, Q => 
                           REGISTERS_39_21_port, QN => n11768);
   REGISTERS_reg_37_21_inst : DFF_X1 port map( D => n13067, CK => n922, Q => 
                           REGISTERS_37_21_port, QN => n11704);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n11883, CK => n922, Q => 
                           REGISTERS_0_21_port, QN => n10478);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n11915, CK => n922, Q => 
                           REGISTERS_1_21_port, QN => n10552);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n11947, CK => n921, Q => 
                           REGISTERS_2_21_port, QN => n10584);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n11979, CK => n921, Q => 
                           REGISTERS_3_21_port, QN => n10616);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n12011, CK => n921, Q => 
                           REGISTERS_4_21_port, QN => n10648);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n12043, CK => n921, Q => 
                           REGISTERS_5_21_port, QN => n10680);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n12075, CK => n921, Q => 
                           REGISTERS_6_21_port, QN => n10712);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n12107, CK => n921, Q => 
                           REGISTERS_7_21_port, QN => n10744);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n12139, CK => n921, Q => 
                           REGISTERS_8_21_port, QN => n10776);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n12171, CK => n921, Q => 
                           REGISTERS_9_21_port, QN => n10808);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n12203, CK => n921, Q => 
                           REGISTERS_10_21_port, QN => n10840);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n12235_port, CK => n921, Q 
                           => REGISTERS_11_21_port, QN => n10872);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n12267_port, CK => n921, Q 
                           => REGISTERS_12_21_port, QN => n10904);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n12299_port, CK => n920, Q 
                           => REGISTERS_13_21_port, QN => n10936);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n12331, CK => n920, Q => 
                           REGISTERS_14_21_port, QN => n10968);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n12363, CK => n920, Q => 
                           REGISTERS_15_21_port, QN => n11000);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n12395, CK => n920, Q => 
                           REGISTERS_16_21_port, QN => n11032);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n12427, CK => n920, Q => 
                           REGISTERS_17_21_port, QN => n11064);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n12459, CK => n920, Q => 
                           REGISTERS_18_21_port, QN => n11096);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n12491, CK => n920, Q => 
                           REGISTERS_19_21_port, QN => n11128);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n12523, CK => n920, Q => 
                           REGISTERS_20_21_port, QN => n11160);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n12555, CK => n920, Q => 
                           REGISTERS_21_21_port, QN => n11192);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n12587, CK => n920, Q => 
                           REGISTERS_22_21_port, QN => n11224);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n12619, CK => n920, Q => 
                           REGISTERS_23_21_port, QN => n11256);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n12651, CK => n919, Q => 
                           REGISTERS_24_21_port, QN => n11288);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n12683, CK => n919, Q => 
                           REGISTERS_25_21_port, QN => n11320);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n12715, CK => n919, Q => 
                           REGISTERS_26_21_port, QN => n11352);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n12747, CK => n919, Q => 
                           REGISTERS_27_21_port, QN => n11384);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n12779, CK => n919, Q => 
                           REGISTERS_28_21_port, QN => n11416);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n12811, CK => n919, Q => 
                           REGISTERS_29_21_port, QN => n11448);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n12843, CK => n919, Q => 
                           REGISTERS_30_21_port, QN => n11480);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n12875, CK => n919, Q => 
                           REGISTERS_31_21_port, QN => n11512);
   REGISTERS_reg_32_21_inst : DFF_X1 port map( D => n12907, CK => n919, Q => 
                           REGISTERS_32_21_port, QN => n11544);
   REGISTERS_reg_33_21_inst : DFF_X1 port map( D => n12939, CK => n919, Q => 
                           REGISTERS_33_21_port, QN => n11576);
   REGISTERS_reg_34_21_inst : DFF_X1 port map( D => n12971, CK => n919, Q => 
                           REGISTERS_34_21_port, QN => n11608);
   REGISTERS_reg_35_21_inst : DFF_X1 port map( D => n13003, CK => n918, Q => 
                           REGISTERS_35_21_port, QN => n11640);
   REGISTERS_reg_36_21_inst : DFF_X1 port map( D => n13035, CK => n922, Q => 
                           REGISTERS_36_21_port, QN => n11672);
   REGISTERS_reg_38_20_inst : DFF_X1 port map( D => n13100, CK => n918, Q => 
                           REGISTERS_38_20_port, QN => n11737);
   REGISTERS_reg_39_20_inst : DFF_X1 port map( D => n13132, CK => n918, Q => 
                           REGISTERS_39_20_port, QN => n11769);
   REGISTERS_reg_37_20_inst : DFF_X1 port map( D => n13068, CK => n918, Q => 
                           REGISTERS_37_20_port, QN => n11705);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n11884, CK => n918, Q => 
                           REGISTERS_0_20_port, QN => n10481);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n11916, CK => n918, Q => 
                           REGISTERS_1_20_port, QN => n10553);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n11948, CK => n918, Q => 
                           REGISTERS_2_20_port, QN => n10585);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n11980, CK => n918, Q => 
                           REGISTERS_3_20_port, QN => n10617);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n12012, CK => n917, Q => 
                           REGISTERS_4_20_port, QN => n10649);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n12044, CK => n917, Q => 
                           REGISTERS_5_20_port, QN => n10681);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n12076, CK => n917, Q => 
                           REGISTERS_6_20_port, QN => n10713);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n12108, CK => n917, Q => 
                           REGISTERS_7_20_port, QN => n10745);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n12140, CK => n917, Q => 
                           REGISTERS_8_20_port, QN => n10777);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n12172, CK => n917, Q => 
                           REGISTERS_9_20_port, QN => n10809);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n12204, CK => n917, Q => 
                           REGISTERS_10_20_port, QN => n10841);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n12236_port, CK => n917, Q 
                           => REGISTERS_11_20_port, QN => n10873);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n12268_port, CK => n917, Q 
                           => REGISTERS_12_20_port, QN => n10905);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n12300_port, CK => n917, Q 
                           => REGISTERS_13_20_port, QN => n10937);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n12332, CK => n917, Q => 
                           REGISTERS_14_20_port, QN => n10969);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n12364, CK => n916, Q => 
                           REGISTERS_15_20_port, QN => n11001);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n12396, CK => n916, Q => 
                           REGISTERS_16_20_port, QN => n11033);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n12428, CK => n916, Q => 
                           REGISTERS_17_20_port, QN => n11065);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n12460, CK => n916, Q => 
                           REGISTERS_18_20_port, QN => n11097);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n12492, CK => n916, Q => 
                           REGISTERS_19_20_port, QN => n11129);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n12524, CK => n916, Q => 
                           REGISTERS_20_20_port, QN => n11161);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n12556, CK => n916, Q => 
                           REGISTERS_21_20_port, QN => n11193);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n12588, CK => n916, Q => 
                           REGISTERS_22_20_port, QN => n11225);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n12620, CK => n916, Q => 
                           REGISTERS_23_20_port, QN => n11257);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n12652, CK => n916, Q => 
                           REGISTERS_24_20_port, QN => n11289);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n12684, CK => n916, Q => 
                           REGISTERS_25_20_port, QN => n11321);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n12716, CK => n915, Q => 
                           REGISTERS_26_20_port, QN => n11353);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n12748, CK => n915, Q => 
                           REGISTERS_27_20_port, QN => n11385);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n12780, CK => n915, Q => 
                           REGISTERS_28_20_port, QN => n11417);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n12812, CK => n915, Q => 
                           REGISTERS_29_20_port, QN => n11449);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n12844, CK => n915, Q => 
                           REGISTERS_30_20_port, QN => n11481);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n12876, CK => n915, Q => 
                           REGISTERS_31_20_port, QN => n11513);
   REGISTERS_reg_32_20_inst : DFF_X1 port map( D => n12908, CK => n915, Q => 
                           REGISTERS_32_20_port, QN => n11545);
   REGISTERS_reg_33_20_inst : DFF_X1 port map( D => n12940, CK => n915, Q => 
                           REGISTERS_33_20_port, QN => n11577);
   REGISTERS_reg_34_20_inst : DFF_X1 port map( D => n12972, CK => n915, Q => 
                           REGISTERS_34_20_port, QN => n11609);
   REGISTERS_reg_35_20_inst : DFF_X1 port map( D => n13004, CK => n915, Q => 
                           REGISTERS_35_20_port, QN => n11641);
   REGISTERS_reg_36_20_inst : DFF_X1 port map( D => n13036, CK => n918, Q => 
                           REGISTERS_36_20_port, QN => n11673);
   REGISTERS_reg_38_19_inst : DFF_X1 port map( D => n13101, CK => n914, Q => 
                           REGISTERS_38_19_port, QN => n11738);
   REGISTERS_reg_39_19_inst : DFF_X1 port map( D => n13133, CK => n914, Q => 
                           REGISTERS_39_19_port, QN => n11770);
   REGISTERS_reg_37_19_inst : DFF_X1 port map( D => n13069, CK => n914, Q => 
                           REGISTERS_37_19_port, QN => n11706);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n11885, CK => n914, Q => 
                           REGISTERS_0_19_port, QN => n10484);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n11917, CK => n914, Q => 
                           REGISTERS_1_19_port, QN => n10554);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n11949, CK => n914, Q => 
                           REGISTERS_2_19_port, QN => n10586);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n11981, CK => n914, Q => 
                           REGISTERS_3_19_port, QN => n10618);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n12013, CK => n914, Q => 
                           REGISTERS_4_19_port, QN => n10650);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n12045, CK => n914, Q => 
                           REGISTERS_5_19_port, QN => n10682);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n12077, CK => n913, Q => 
                           REGISTERS_6_19_port, QN => n10714);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n12109, CK => n913, Q => 
                           REGISTERS_7_19_port, QN => n10746);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n12141, CK => n913, Q => 
                           REGISTERS_8_19_port, QN => n10778);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n12173, CK => n913, Q => 
                           REGISTERS_9_19_port, QN => n10810);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n12205_port, CK => n913, Q 
                           => REGISTERS_10_19_port, QN => n10842);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n12237_port, CK => n913, Q 
                           => REGISTERS_11_19_port, QN => n10874);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n12269_port, CK => n913, Q 
                           => REGISTERS_12_19_port, QN => n10906);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n12301, CK => n913, Q => 
                           REGISTERS_13_19_port, QN => n10938);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n12333, CK => n913, Q => 
                           REGISTERS_14_19_port, QN => n10970);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n12365, CK => n913, Q => 
                           REGISTERS_15_19_port, QN => n11002);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n12397, CK => n913, Q => 
                           REGISTERS_16_19_port, QN => n11034);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n12429, CK => n912, Q => 
                           REGISTERS_17_19_port, QN => n11066);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n12461, CK => n912, Q => 
                           REGISTERS_18_19_port, QN => n11098);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n12493, CK => n912, Q => 
                           REGISTERS_19_19_port, QN => n11130);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n12525, CK => n912, Q => 
                           REGISTERS_20_19_port, QN => n11162);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n12557, CK => n912, Q => 
                           REGISTERS_21_19_port, QN => n11194);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n12589, CK => n912, Q => 
                           REGISTERS_22_19_port, QN => n11226);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n12621, CK => n912, Q => 
                           REGISTERS_23_19_port, QN => n11258);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n12653, CK => n912, Q => 
                           REGISTERS_24_19_port, QN => n11290);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n12685, CK => n912, Q => 
                           REGISTERS_25_19_port, QN => n11322);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n12717, CK => n912, Q => 
                           REGISTERS_26_19_port, QN => n11354);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n12749, CK => n912, Q => 
                           REGISTERS_27_19_port, QN => n11386);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n12781, CK => n911, Q => 
                           REGISTERS_28_19_port, QN => n11418);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n12813, CK => n911, Q => 
                           REGISTERS_29_19_port, QN => n11450);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n12845, CK => n911, Q => 
                           REGISTERS_30_19_port, QN => n11482);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n12877, CK => n911, Q => 
                           REGISTERS_31_19_port, QN => n11514);
   REGISTERS_reg_32_19_inst : DFF_X1 port map( D => n12909, CK => n911, Q => 
                           REGISTERS_32_19_port, QN => n11546);
   REGISTERS_reg_33_19_inst : DFF_X1 port map( D => n12941, CK => n911, Q => 
                           REGISTERS_33_19_port, QN => n11578);
   REGISTERS_reg_34_19_inst : DFF_X1 port map( D => n12973, CK => n911, Q => 
                           REGISTERS_34_19_port, QN => n11610);
   REGISTERS_reg_35_19_inst : DFF_X1 port map( D => n13005, CK => n911, Q => 
                           REGISTERS_35_19_port, QN => n11642);
   REGISTERS_reg_36_19_inst : DFF_X1 port map( D => n13037, CK => n914, Q => 
                           REGISTERS_36_19_port, QN => n11674);
   REGISTERS_reg_38_18_inst : DFF_X1 port map( D => n13102, CK => n910, Q => 
                           REGISTERS_38_18_port, QN => n11739);
   REGISTERS_reg_39_18_inst : DFF_X1 port map( D => n13134, CK => n910, Q => 
                           REGISTERS_39_18_port, QN => n11771);
   REGISTERS_reg_37_18_inst : DFF_X1 port map( D => n13070, CK => n910, Q => 
                           REGISTERS_37_18_port, QN => n11707);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n11886, CK => n910, Q => 
                           REGISTERS_0_18_port, QN => n10487);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n11918, CK => n910, Q => 
                           REGISTERS_1_18_port, QN => n10555);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n11950, CK => n910, Q => 
                           REGISTERS_2_18_port, QN => n10587);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n11982, CK => n910, Q => 
                           REGISTERS_3_18_port, QN => n10619);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n12014, CK => n910, Q => 
                           REGISTERS_4_18_port, QN => n10651);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n12046, CK => n910, Q => 
                           REGISTERS_5_18_port, QN => n10683);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n12078, CK => n910, Q => 
                           REGISTERS_6_18_port, QN => n10715);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n12110, CK => n910, Q => 
                           REGISTERS_7_18_port, QN => n10747);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n12142, CK => n909, Q => 
                           REGISTERS_8_18_port, QN => n10779);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n12174, CK => n909, Q => 
                           REGISTERS_9_18_port, QN => n10811);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n12206_port, CK => n909, Q 
                           => REGISTERS_10_18_port, QN => n10843);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n12238_port, CK => n909, Q 
                           => REGISTERS_11_18_port, QN => n10875);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n12270_port, CK => n909, Q 
                           => REGISTERS_12_18_port, QN => n10907);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n12302, CK => n909, Q => 
                           REGISTERS_13_18_port, QN => n10939);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n12334, CK => n909, Q => 
                           REGISTERS_14_18_port, QN => n10971);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n12366, CK => n909, Q => 
                           REGISTERS_15_18_port, QN => n11003);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n12398, CK => n909, Q => 
                           REGISTERS_16_18_port, QN => n11035);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n12430, CK => n909, Q => 
                           REGISTERS_17_18_port, QN => n11067);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n12462, CK => n909, Q => 
                           REGISTERS_18_18_port, QN => n11099);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n12494, CK => n908, Q => 
                           REGISTERS_19_18_port, QN => n11131);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n12526, CK => n908, Q => 
                           REGISTERS_20_18_port, QN => n11163);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n12558, CK => n908, Q => 
                           REGISTERS_21_18_port, QN => n11195);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n12590, CK => n908, Q => 
                           REGISTERS_22_18_port, QN => n11227);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n12622, CK => n908, Q => 
                           REGISTERS_23_18_port, QN => n11259);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n12654, CK => n908, Q => 
                           REGISTERS_24_18_port, QN => n11291);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n12686, CK => n908, Q => 
                           REGISTERS_25_18_port, QN => n11323);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n12718, CK => n908, Q => 
                           REGISTERS_26_18_port, QN => n11355);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n12750, CK => n908, Q => 
                           REGISTERS_27_18_port, QN => n11387);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n12782, CK => n908, Q => 
                           REGISTERS_28_18_port, QN => n11419);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n12814, CK => n908, Q => 
                           REGISTERS_29_18_port, QN => n11451);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n12846, CK => n907, Q => 
                           REGISTERS_30_18_port, QN => n11483);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n12878, CK => n907, Q => 
                           REGISTERS_31_18_port, QN => n11515);
   REGISTERS_reg_32_18_inst : DFF_X1 port map( D => n12910, CK => n907, Q => 
                           REGISTERS_32_18_port, QN => n11547);
   REGISTERS_reg_33_18_inst : DFF_X1 port map( D => n12942, CK => n907, Q => 
                           REGISTERS_33_18_port, QN => n11579);
   REGISTERS_reg_34_18_inst : DFF_X1 port map( D => n12974, CK => n907, Q => 
                           REGISTERS_34_18_port, QN => n11611);
   REGISTERS_reg_35_18_inst : DFF_X1 port map( D => n13006, CK => n907, Q => 
                           REGISTERS_35_18_port, QN => n11643);
   REGISTERS_reg_36_18_inst : DFF_X1 port map( D => n13038, CK => n911, Q => 
                           REGISTERS_36_18_port, QN => n11675);
   REGISTERS_reg_38_17_inst : DFF_X1 port map( D => n13103, CK => n907, Q => 
                           REGISTERS_38_17_port, QN => n11740);
   REGISTERS_reg_39_17_inst : DFF_X1 port map( D => n13135, CK => n907, Q => 
                           REGISTERS_39_17_port, QN => n11772);
   REGISTERS_reg_37_17_inst : DFF_X1 port map( D => n13071, CK => n906, Q => 
                           REGISTERS_37_17_port, QN => n11708);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n11887, CK => n906, Q => 
                           REGISTERS_0_17_port, QN => n10490);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n11919, CK => n906, Q => 
                           REGISTERS_1_17_port, QN => n10556);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n11951, CK => n906, Q => 
                           REGISTERS_2_17_port, QN => n10588);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n11983, CK => n906, Q => 
                           REGISTERS_3_17_port, QN => n10620);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n12015, CK => n906, Q => 
                           REGISTERS_4_17_port, QN => n10652);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n12047, CK => n906, Q => 
                           REGISTERS_5_17_port, QN => n10684);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n12079, CK => n906, Q => 
                           REGISTERS_6_17_port, QN => n10716);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n12111, CK => n906, Q => 
                           REGISTERS_7_17_port, QN => n10748);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n12143, CK => n906, Q => 
                           REGISTERS_8_17_port, QN => n10780);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n12175, CK => n906, Q => 
                           REGISTERS_9_17_port, QN => n10812);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n12207_port, CK => n905, Q 
                           => REGISTERS_10_17_port, QN => n10844);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n12239_port, CK => n905, Q 
                           => REGISTERS_11_17_port, QN => n10876);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n12271_port, CK => n905, Q 
                           => REGISTERS_12_17_port, QN => n10908);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n12303, CK => n905, Q => 
                           REGISTERS_13_17_port, QN => n10940);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n12335, CK => n905, Q => 
                           REGISTERS_14_17_port, QN => n10972);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n12367, CK => n905, Q => 
                           REGISTERS_15_17_port, QN => n11004);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n12399, CK => n905, Q => 
                           REGISTERS_16_17_port, QN => n11036);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n12431, CK => n905, Q => 
                           REGISTERS_17_17_port, QN => n11068);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n12463, CK => n905, Q => 
                           REGISTERS_18_17_port, QN => n11100);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n12495, CK => n905, Q => 
                           REGISTERS_19_17_port, QN => n11132);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n12527, CK => n905, Q => 
                           REGISTERS_20_17_port, QN => n11164);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n12559, CK => n904, Q => 
                           REGISTERS_21_17_port, QN => n11196);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n12591, CK => n904, Q => 
                           REGISTERS_22_17_port, QN => n11228);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n12623, CK => n904, Q => 
                           REGISTERS_23_17_port, QN => n11260);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n12655, CK => n904, Q => 
                           REGISTERS_24_17_port, QN => n11292);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n12687, CK => n904, Q => 
                           REGISTERS_25_17_port, QN => n11324);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n12719, CK => n904, Q => 
                           REGISTERS_26_17_port, QN => n11356);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n12751, CK => n904, Q => 
                           REGISTERS_27_17_port, QN => n11388);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n12783, CK => n904, Q => 
                           REGISTERS_28_17_port, QN => n11420);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n12815, CK => n904, Q => 
                           REGISTERS_29_17_port, QN => n11452);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n12847, CK => n904, Q => 
                           REGISTERS_30_17_port, QN => n11484);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n12879, CK => n904, Q => 
                           REGISTERS_31_17_port, QN => n11516);
   REGISTERS_reg_32_17_inst : DFF_X1 port map( D => n12911, CK => n903, Q => 
                           REGISTERS_32_17_port, QN => n11548);
   REGISTERS_reg_33_17_inst : DFF_X1 port map( D => n12943, CK => n903, Q => 
                           REGISTERS_33_17_port, QN => n11580);
   REGISTERS_reg_34_17_inst : DFF_X1 port map( D => n12975, CK => n903, Q => 
                           REGISTERS_34_17_port, QN => n11612);
   REGISTERS_reg_35_17_inst : DFF_X1 port map( D => n13007, CK => n903, Q => 
                           REGISTERS_35_17_port, QN => n11644);
   REGISTERS_reg_36_17_inst : DFF_X1 port map( D => n13039, CK => n907, Q => 
                           REGISTERS_36_17_port, QN => n11676);
   REGISTERS_reg_38_16_inst : DFF_X1 port map( D => n13104, CK => n964, Q => 
                           REGISTERS_38_16_port, QN => n11741);
   REGISTERS_reg_39_16_inst : DFF_X1 port map( D => n13136, CK => n964, Q => 
                           REGISTERS_39_16_port, QN => n11773);
   REGISTERS_reg_37_16_inst : DFF_X1 port map( D => n13072, CK => n964, Q => 
                           REGISTERS_37_16_port, QN => n11709);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n11888, CK => n964, Q => 
                           REGISTERS_0_16_port, QN => n10493);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n11920, CK => n964, Q => 
                           REGISTERS_1_16_port, QN => n10557);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n11952, CK => n963, Q => 
                           REGISTERS_2_16_port, QN => n10589);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n11984, CK => n963, Q => 
                           REGISTERS_3_16_port, QN => n10621);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n12016, CK => n963, Q => 
                           REGISTERS_4_16_port, QN => n10653);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n12048, CK => n963, Q => 
                           REGISTERS_5_16_port, QN => n10685);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n12080, CK => n963, Q => 
                           REGISTERS_6_16_port, QN => n10717);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n12112, CK => n963, Q => 
                           REGISTERS_7_16_port, QN => n10749);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n12144, CK => n963, Q => 
                           REGISTERS_8_16_port, QN => n10781);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n12176, CK => n963, Q => 
                           REGISTERS_9_16_port, QN => n10813);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n12208_port, CK => n963, Q 
                           => REGISTERS_10_16_port, QN => n10845);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n12240_port, CK => n963, Q 
                           => REGISTERS_11_16_port, QN => n10877);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n12272_port, CK => n963, Q 
                           => REGISTERS_12_16_port, QN => n10909);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n12304, CK => n962, Q => 
                           REGISTERS_13_16_port, QN => n10941);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n12336, CK => n962, Q => 
                           REGISTERS_14_16_port, QN => n10973);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n12368, CK => n962, Q => 
                           REGISTERS_15_16_port, QN => n11005);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n12400, CK => n962, Q => 
                           REGISTERS_16_16_port, QN => n11037);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n12432, CK => n962, Q => 
                           REGISTERS_17_16_port, QN => n11069);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n12464, CK => n962, Q => 
                           REGISTERS_18_16_port, QN => n11101);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n12496, CK => n962, Q => 
                           REGISTERS_19_16_port, QN => n11133);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n12528, CK => n962, Q => 
                           REGISTERS_20_16_port, QN => n11165);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n12560, CK => n962, Q => 
                           REGISTERS_21_16_port, QN => n11197);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n12592, CK => n962, Q => 
                           REGISTERS_22_16_port, QN => n11229);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n12624, CK => n962, Q => 
                           REGISTERS_23_16_port, QN => n11261);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n12656, CK => n961, Q => 
                           REGISTERS_24_16_port, QN => n11293);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n12688, CK => n961, Q => 
                           REGISTERS_25_16_port, QN => n11325);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n12720, CK => n961, Q => 
                           REGISTERS_26_16_port, QN => n11357);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n12752, CK => n961, Q => 
                           REGISTERS_27_16_port, QN => n11389);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n12784, CK => n961, Q => 
                           REGISTERS_28_16_port, QN => n11421);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n12816, CK => n961, Q => 
                           REGISTERS_29_16_port, QN => n11453);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n12848, CK => n961, Q => 
                           REGISTERS_30_16_port, QN => n11485);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n12880, CK => n961, Q => 
                           REGISTERS_31_16_port, QN => n11517);
   REGISTERS_reg_32_16_inst : DFF_X1 port map( D => n12912, CK => n961, Q => 
                           REGISTERS_32_16_port, QN => n11549);
   REGISTERS_reg_33_16_inst : DFF_X1 port map( D => n12944, CK => n961, Q => 
                           REGISTERS_33_16_port, QN => n11581);
   REGISTERS_reg_34_16_inst : DFF_X1 port map( D => n12976, CK => n961, Q => 
                           REGISTERS_34_16_port, QN => n11613);
   REGISTERS_reg_35_16_inst : DFF_X1 port map( D => n13008, CK => n960, Q => 
                           REGISTERS_35_16_port, QN => n11645);
   REGISTERS_reg_36_16_inst : DFF_X1 port map( D => n13040, CK => n964, Q => 
                           REGISTERS_36_16_port, QN => n11677);
   REGISTERS_reg_38_15_inst : DFF_X1 port map( D => n13105, CK => n903, Q => 
                           REGISTERS_38_15_port, QN => n11742);
   REGISTERS_reg_39_15_inst : DFF_X1 port map( D => n13137, CK => n903, Q => 
                           REGISTERS_39_15_port, QN => n11774);
   REGISTERS_reg_37_15_inst : DFF_X1 port map( D => n13073, CK => n903, Q => 
                           REGISTERS_37_15_port, QN => n11710);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n11889, CK => n903, Q => 
                           REGISTERS_0_15_port, QN => n10496);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n11921, CK => n902, Q => 
                           REGISTERS_1_15_port, QN => n10558);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n11953, CK => n902, Q => 
                           REGISTERS_2_15_port, QN => n10590);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n11985, CK => n902, Q => 
                           REGISTERS_3_15_port, QN => n10622);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n12017, CK => n902, Q => 
                           REGISTERS_4_15_port, QN => n10654);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n12049, CK => n902, Q => 
                           REGISTERS_5_15_port, QN => n10686);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n12081, CK => n902, Q => 
                           REGISTERS_6_15_port, QN => n10718);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n12113, CK => n902, Q => 
                           REGISTERS_7_15_port, QN => n10750);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n12145, CK => n902, Q => 
                           REGISTERS_8_15_port, QN => n10782);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n12177, CK => n902, Q => 
                           REGISTERS_9_15_port, QN => n10814);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n12209_port, CK => n902, Q 
                           => REGISTERS_10_15_port, QN => n10846);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n12241_port, CK => n902, Q 
                           => REGISTERS_11_15_port, QN => n10878);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n12273_port, CK => n901, Q 
                           => REGISTERS_12_15_port, QN => n10910);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n12305, CK => n901, Q => 
                           REGISTERS_13_15_port, QN => n10942);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n12337, CK => n901, Q => 
                           REGISTERS_14_15_port, QN => n10974);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n12369, CK => n901, Q => 
                           REGISTERS_15_15_port, QN => n11006);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n12401, CK => n901, Q => 
                           REGISTERS_16_15_port, QN => n11038);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n12433, CK => n901, Q => 
                           REGISTERS_17_15_port, QN => n11070);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n12465, CK => n901, Q => 
                           REGISTERS_18_15_port, QN => n11102);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n12497, CK => n901, Q => 
                           REGISTERS_19_15_port, QN => n11134);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n12529, CK => n901, Q => 
                           REGISTERS_20_15_port, QN => n11166);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n12561, CK => n901, Q => 
                           REGISTERS_21_15_port, QN => n11198);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n12593, CK => n901, Q => 
                           REGISTERS_22_15_port, QN => n11230);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n12625, CK => n900, Q => 
                           REGISTERS_23_15_port, QN => n11262);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n12657, CK => n900, Q => 
                           REGISTERS_24_15_port, QN => n11294);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n12689, CK => n900, Q => 
                           REGISTERS_25_15_port, QN => n11326);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n12721, CK => n900, Q => 
                           REGISTERS_26_15_port, QN => n11358);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n12753, CK => n900, Q => 
                           REGISTERS_27_15_port, QN => n11390);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n12785, CK => n900, Q => 
                           REGISTERS_28_15_port, QN => n11422);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n12817, CK => n900, Q => 
                           REGISTERS_29_15_port, QN => n11454);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n12849, CK => n900, Q => 
                           REGISTERS_30_15_port, QN => n11486);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n12881, CK => n900, Q => 
                           REGISTERS_31_15_port, QN => n11518);
   REGISTERS_reg_32_15_inst : DFF_X1 port map( D => n12913, CK => n900, Q => 
                           REGISTERS_32_15_port, QN => n11550);
   REGISTERS_reg_33_15_inst : DFF_X1 port map( D => n12945, CK => n900, Q => 
                           REGISTERS_33_15_port, QN => n11582);
   REGISTERS_reg_34_15_inst : DFF_X1 port map( D => n12977, CK => n899, Q => 
                           REGISTERS_34_15_port, QN => n11614);
   REGISTERS_reg_35_15_inst : DFF_X1 port map( D => n13009, CK => n899, Q => 
                           REGISTERS_35_15_port, QN => n11646);
   REGISTERS_reg_36_15_inst : DFF_X1 port map( D => n13041, CK => n903, Q => 
                           REGISTERS_36_15_port, QN => n11678);
   REGISTERS_reg_38_14_inst : DFF_X1 port map( D => n13106, CK => n880, Q => 
                           REGISTERS_38_14_port, QN => n11743);
   REGISTERS_reg_39_14_inst : DFF_X1 port map( D => n13138, CK => n880, Q => 
                           REGISTERS_39_14_port, QN => n11775);
   REGISTERS_reg_37_14_inst : DFF_X1 port map( D => n13074, CK => n880, Q => 
                           REGISTERS_37_14_port, QN => n11711);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n11890, CK => n880, Q => 
                           REGISTERS_0_14_port, QN => n10499);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n11922, CK => n880, Q => 
                           REGISTERS_1_14_port, QN => n10559);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n11954, CK => n879, Q => 
                           REGISTERS_2_14_port, QN => n10591);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n11986, CK => n879, Q => 
                           REGISTERS_3_14_port, QN => n10623);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n12018, CK => n879, Q => 
                           REGISTERS_4_14_port, QN => n10655);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n12050, CK => n879, Q => 
                           REGISTERS_5_14_port, QN => n10687);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n12082, CK => n879, Q => 
                           REGISTERS_6_14_port, QN => n10719);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n12114, CK => n879, Q => 
                           REGISTERS_7_14_port, QN => n10751);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n12146, CK => n879, Q => 
                           REGISTERS_8_14_port, QN => n10783);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n12178, CK => n879, Q => 
                           REGISTERS_9_14_port, QN => n10815);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n12210_port, CK => n879, Q 
                           => REGISTERS_10_14_port, QN => n10847);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n12242_port, CK => n879, Q 
                           => REGISTERS_11_14_port, QN => n10879);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n12274_port, CK => n879, Q 
                           => REGISTERS_12_14_port, QN => n10911);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n12306, CK => n878, Q => 
                           REGISTERS_13_14_port, QN => n10943);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n12338, CK => n878, Q => 
                           REGISTERS_14_14_port, QN => n10975);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n12370, CK => n878, Q => 
                           REGISTERS_15_14_port, QN => n11007);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n12402, CK => n878, Q => 
                           REGISTERS_16_14_port, QN => n11039);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n12434, CK => n878, Q => 
                           REGISTERS_17_14_port, QN => n11071);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n12466, CK => n878, Q => 
                           REGISTERS_18_14_port, QN => n11103);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n12498, CK => n878, Q => 
                           REGISTERS_19_14_port, QN => n11135);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n12530, CK => n878, Q => 
                           REGISTERS_20_14_port, QN => n11167);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n12562, CK => n878, Q => 
                           REGISTERS_21_14_port, QN => n11199);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n12594, CK => n878, Q => 
                           REGISTERS_22_14_port, QN => n11231);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n12626, CK => n878, Q => 
                           REGISTERS_23_14_port, QN => n11263);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n12658, CK => n877, Q => 
                           REGISTERS_24_14_port, QN => n11295);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n12690, CK => n877, Q => 
                           REGISTERS_25_14_port, QN => n11327);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n12722, CK => n877, Q => 
                           REGISTERS_26_14_port, QN => n11359);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n12754, CK => n877, Q => 
                           REGISTERS_27_14_port, QN => n11391);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n12786, CK => n877, Q => 
                           REGISTERS_28_14_port, QN => n11423);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n12818, CK => n877, Q => 
                           REGISTERS_29_14_port, QN => n11455);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n12850, CK => n877, Q => 
                           REGISTERS_30_14_port, QN => n11487);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n12882, CK => n877, Q => 
                           REGISTERS_31_14_port, QN => n11519);
   REGISTERS_reg_32_14_inst : DFF_X1 port map( D => n12914, CK => n877, Q => 
                           REGISTERS_32_14_port, QN => n11551);
   REGISTERS_reg_33_14_inst : DFF_X1 port map( D => n12946, CK => n877, Q => 
                           REGISTERS_33_14_port, QN => n11583);
   REGISTERS_reg_34_14_inst : DFF_X1 port map( D => n12978, CK => n877, Q => 
                           REGISTERS_34_14_port, QN => n11615);
   REGISTERS_reg_35_14_inst : DFF_X1 port map( D => n13010, CK => n876, Q => 
                           REGISTERS_35_14_port, QN => n11647);
   REGISTERS_reg_36_14_inst : DFF_X1 port map( D => n13042, CK => n880, Q => 
                           REGISTERS_36_14_port, QN => n11679);
   REGISTERS_reg_38_13_inst : DFF_X1 port map( D => n13107, CK => n876, Q => 
                           REGISTERS_38_13_port, QN => n11744);
   REGISTERS_reg_39_13_inst : DFF_X1 port map( D => n13139, CK => n876, Q => 
                           REGISTERS_39_13_port, QN => n11776);
   REGISTERS_reg_37_13_inst : DFF_X1 port map( D => n13075, CK => n876, Q => 
                           REGISTERS_37_13_port, QN => n11712);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n11891, CK => n876, Q => 
                           REGISTERS_0_13_port, QN => n10502);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n11923, CK => n876, Q => 
                           REGISTERS_1_13_port, QN => n10560);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n11955, CK => n876, Q => 
                           REGISTERS_2_13_port, QN => n10592);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n11987, CK => n876, Q => 
                           REGISTERS_3_13_port, QN => n10624);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n12019, CK => n875, Q => 
                           REGISTERS_4_13_port, QN => n10656);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n12051, CK => n875, Q => 
                           REGISTERS_5_13_port, QN => n10688);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n12083, CK => n875, Q => 
                           REGISTERS_6_13_port, QN => n10720);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n12115, CK => n875, Q => 
                           REGISTERS_7_13_port, QN => n10752);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n12147, CK => n875, Q => 
                           REGISTERS_8_13_port, QN => n10784);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n12179, CK => n875, Q => 
                           REGISTERS_9_13_port, QN => n10816);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n12211_port, CK => n875, Q 
                           => REGISTERS_10_13_port, QN => n10848);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n12243_port, CK => n875, Q 
                           => REGISTERS_11_13_port, QN => n10880);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n12275_port, CK => n875, Q 
                           => REGISTERS_12_13_port, QN => n10912);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n12307, CK => n875, Q => 
                           REGISTERS_13_13_port, QN => n10944);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n12339, CK => n875, Q => 
                           REGISTERS_14_13_port, QN => n10976);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n12371, CK => n874, Q => 
                           REGISTERS_15_13_port, QN => n11008);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n12403, CK => n874, Q => 
                           REGISTERS_16_13_port, QN => n11040);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n12435, CK => n874, Q => 
                           REGISTERS_17_13_port, QN => n11072);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n12467, CK => n874, Q => 
                           REGISTERS_18_13_port, QN => n11104);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n12499, CK => n874, Q => 
                           REGISTERS_19_13_port, QN => n11136);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n12531, CK => n874, Q => 
                           REGISTERS_20_13_port, QN => n11168);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n12563, CK => n874, Q => 
                           REGISTERS_21_13_port, QN => n11200);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n12595, CK => n874, Q => 
                           REGISTERS_22_13_port, QN => n11232);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n12627, CK => n874, Q => 
                           REGISTERS_23_13_port, QN => n11264);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n12659, CK => n874, Q => 
                           REGISTERS_24_13_port, QN => n11296);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n12691, CK => n874, Q => 
                           REGISTERS_25_13_port, QN => n11328);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n12723, CK => n873, Q => 
                           REGISTERS_26_13_port, QN => n11360);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n12755, CK => n873, Q => 
                           REGISTERS_27_13_port, QN => n11392);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n12787, CK => n873, Q => 
                           REGISTERS_28_13_port, QN => n11424);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n12819, CK => n873, Q => 
                           REGISTERS_29_13_port, QN => n11456);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n12851, CK => n873, Q => 
                           REGISTERS_30_13_port, QN => n11488);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n12883, CK => n873, Q => 
                           REGISTERS_31_13_port, QN => n11520);
   REGISTERS_reg_32_13_inst : DFF_X1 port map( D => n12915, CK => n873, Q => 
                           REGISTERS_32_13_port, QN => n11552);
   REGISTERS_reg_33_13_inst : DFF_X1 port map( D => n12947, CK => n873, Q => 
                           REGISTERS_33_13_port, QN => n11584);
   REGISTERS_reg_34_13_inst : DFF_X1 port map( D => n12979, CK => n873, Q => 
                           REGISTERS_34_13_port, QN => n11616);
   REGISTERS_reg_35_13_inst : DFF_X1 port map( D => n13011, CK => n873, Q => 
                           REGISTERS_35_13_port, QN => n11648);
   REGISTERS_reg_36_13_inst : DFF_X1 port map( D => n13043, CK => n876, Q => 
                           REGISTERS_36_13_port, QN => n11680);
   REGISTERS_reg_38_12_inst : DFF_X1 port map( D => n13108, CK => n949, Q => 
                           REGISTERS_38_12_port, QN => n11745);
   REGISTERS_reg_39_12_inst : DFF_X1 port map( D => n13140, CK => n949, Q => 
                           REGISTERS_39_12_port, QN => n11777);
   REGISTERS_reg_37_12_inst : DFF_X1 port map( D => n13076, CK => n948, Q => 
                           REGISTERS_37_12_port, QN => n11713);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n11892, CK => n948, Q => 
                           REGISTERS_0_12_port, QN => n10505);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n11924, CK => n948, Q => 
                           REGISTERS_1_12_port, QN => n10561);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n11956, CK => n948, Q => 
                           REGISTERS_2_12_port, QN => n10593);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n11988, CK => n948, Q => 
                           REGISTERS_3_12_port, QN => n10625);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n12020, CK => n948, Q => 
                           REGISTERS_4_12_port, QN => n10657);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n12052, CK => n948, Q => 
                           REGISTERS_5_12_port, QN => n10689);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n12084, CK => n948, Q => 
                           REGISTERS_6_12_port, QN => n10721);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n12116, CK => n948, Q => 
                           REGISTERS_7_12_port, QN => n10753);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n12148, CK => n948, Q => 
                           REGISTERS_8_12_port, QN => n10785);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n12180, CK => n948, Q => 
                           REGISTERS_9_12_port, QN => n10817);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n12212_port, CK => n947, Q 
                           => REGISTERS_10_12_port, QN => n10849);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n12244_port, CK => n947, Q 
                           => REGISTERS_11_12_port, QN => n10881);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n12276_port, CK => n947, Q 
                           => REGISTERS_12_12_port, QN => n10913);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n12308, CK => n947, Q => 
                           REGISTERS_13_12_port, QN => n10945);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n12340, CK => n947, Q => 
                           REGISTERS_14_12_port, QN => n10977);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n12372, CK => n947, Q => 
                           REGISTERS_15_12_port, QN => n11009);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n12404, CK => n947, Q => 
                           REGISTERS_16_12_port, QN => n11041);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n12436, CK => n947, Q => 
                           REGISTERS_17_12_port, QN => n11073);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n12468, CK => n947, Q => 
                           REGISTERS_18_12_port, QN => n11105);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n12500, CK => n947, Q => 
                           REGISTERS_19_12_port, QN => n11137);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n12532, CK => n947, Q => 
                           REGISTERS_20_12_port, QN => n11169);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n12564, CK => n946, Q => 
                           REGISTERS_21_12_port, QN => n11201);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n12596, CK => n946, Q => 
                           REGISTERS_22_12_port, QN => n11233);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n12628, CK => n946, Q => 
                           REGISTERS_23_12_port, QN => n11265);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n12660, CK => n946, Q => 
                           REGISTERS_24_12_port, QN => n11297);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n12692, CK => n946, Q => 
                           REGISTERS_25_12_port, QN => n11329);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n12724, CK => n946, Q => 
                           REGISTERS_26_12_port, QN => n11361);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n12756, CK => n946, Q => 
                           REGISTERS_27_12_port, QN => n11393);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n12788, CK => n946, Q => 
                           REGISTERS_28_12_port, QN => n11425);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n12820, CK => n946, Q => 
                           REGISTERS_29_12_port, QN => n11457);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n12852, CK => n946, Q => 
                           REGISTERS_30_12_port, QN => n11489);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n12884, CK => n946, Q => 
                           REGISTERS_31_12_port, QN => n11521);
   REGISTERS_reg_32_12_inst : DFF_X1 port map( D => n12916, CK => n945, Q => 
                           REGISTERS_32_12_port, QN => n11553);
   REGISTERS_reg_33_12_inst : DFF_X1 port map( D => n12948, CK => n945, Q => 
                           REGISTERS_33_12_port, QN => n11585);
   REGISTERS_reg_34_12_inst : DFF_X1 port map( D => n12980, CK => n945, Q => 
                           REGISTERS_34_12_port, QN => n11617);
   REGISTERS_reg_35_12_inst : DFF_X1 port map( D => n13012, CK => n945, Q => 
                           REGISTERS_35_12_port, QN => n11649);
   REGISTERS_reg_36_12_inst : DFF_X1 port map( D => n13044, CK => n949, Q => 
                           REGISTERS_36_12_port, QN => n11681);
   REGISTERS_reg_38_11_inst : DFF_X1 port map( D => n13109, CK => n884, Q => 
                           REGISTERS_38_11_port, QN => n11746);
   REGISTERS_reg_39_11_inst : DFF_X1 port map( D => n13141, CK => n884, Q => 
                           REGISTERS_39_11_port, QN => n11778);
   REGISTERS_reg_37_11_inst : DFF_X1 port map( D => n13077, CK => n884, Q => 
                           REGISTERS_37_11_port, QN => n11714);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n11893, CK => n883, Q => 
                           REGISTERS_0_11_port, QN => n10508);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n11925, CK => n883, Q => 
                           REGISTERS_1_11_port, QN => n10562);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n11957, CK => n883, Q => 
                           REGISTERS_2_11_port, QN => n10594);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n11989, CK => n883, Q => 
                           REGISTERS_3_11_port, QN => n10626);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n12021, CK => n883, Q => 
                           REGISTERS_4_11_port, QN => n10658);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n12053, CK => n883, Q => 
                           REGISTERS_5_11_port, QN => n10690);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n12085, CK => n883, Q => 
                           REGISTERS_6_11_port, QN => n10722);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n12117, CK => n883, Q => 
                           REGISTERS_7_11_port, QN => n10754);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n12149, CK => n883, Q => 
                           REGISTERS_8_11_port, QN => n10786);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n12181, CK => n883, Q => 
                           REGISTERS_9_11_port, QN => n10818);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n12213_port, CK => n883, Q 
                           => REGISTERS_10_11_port, QN => n10850);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n12245_port, CK => n882, Q 
                           => REGISTERS_11_11_port, QN => n10882);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n12277_port, CK => n882, Q 
                           => REGISTERS_12_11_port, QN => n10914);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n12309, CK => n882, Q => 
                           REGISTERS_13_11_port, QN => n10946);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n12341, CK => n882, Q => 
                           REGISTERS_14_11_port, QN => n10978);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n12373, CK => n882, Q => 
                           REGISTERS_15_11_port, QN => n11010);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n12405, CK => n882, Q => 
                           REGISTERS_16_11_port, QN => n11042);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n12437, CK => n882, Q => 
                           REGISTERS_17_11_port, QN => n11074);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n12469, CK => n882, Q => 
                           REGISTERS_18_11_port, QN => n11106);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n12501, CK => n882, Q => 
                           REGISTERS_19_11_port, QN => n11138);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n12533, CK => n882, Q => 
                           REGISTERS_20_11_port, QN => n11170);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n12565, CK => n882, Q => 
                           REGISTERS_21_11_port, QN => n11202);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n12597, CK => n881, Q => 
                           REGISTERS_22_11_port, QN => n11234);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n12629, CK => n881, Q => 
                           REGISTERS_23_11_port, QN => n11266);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n12661, CK => n881, Q => 
                           REGISTERS_24_11_port, QN => n11298);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n12693, CK => n881, Q => 
                           REGISTERS_25_11_port, QN => n11330);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n12725, CK => n881, Q => 
                           REGISTERS_26_11_port, QN => n11362);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n12757, CK => n881, Q => 
                           REGISTERS_27_11_port, QN => n11394);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n12789, CK => n881, Q => 
                           REGISTERS_28_11_port, QN => n11426);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n12821, CK => n881, Q => 
                           REGISTERS_29_11_port, QN => n11458);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n12853, CK => n881, Q => 
                           REGISTERS_30_11_port, QN => n11490);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n12885, CK => n881, Q => 
                           REGISTERS_31_11_port, QN => n11522);
   REGISTERS_reg_32_11_inst : DFF_X1 port map( D => n12917, CK => n881, Q => 
                           REGISTERS_32_11_port, QN => n11554);
   REGISTERS_reg_33_11_inst : DFF_X1 port map( D => n12949, CK => n880, Q => 
                           REGISTERS_33_11_port, QN => n11586);
   REGISTERS_reg_34_11_inst : DFF_X1 port map( D => n12981, CK => n880, Q => 
                           REGISTERS_34_11_port, QN => n11618);
   REGISTERS_reg_35_11_inst : DFF_X1 port map( D => n13013, CK => n880, Q => 
                           REGISTERS_35_11_port, QN => n11650);
   REGISTERS_reg_36_11_inst : DFF_X1 port map( D => n13045, CK => n884, Q => 
                           REGISTERS_36_11_port, QN => n11682);
   REGISTERS_reg_38_10_inst : DFF_X1 port map( D => n13110, CK => n872, Q => 
                           REGISTERS_38_10_port, QN => n11747);
   REGISTERS_reg_39_10_inst : DFF_X1 port map( D => n13142, CK => n872, Q => 
                           REGISTERS_39_10_port, QN => n11779);
   REGISTERS_reg_37_10_inst : DFF_X1 port map( D => n13078, CK => n872, Q => 
                           REGISTERS_37_10_port, QN => n11715);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n11894, CK => n872, Q => 
                           REGISTERS_0_10_port, QN => n10511);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n11926, CK => n872, Q => 
                           REGISTERS_1_10_port, QN => n10563);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n11958, CK => n872, Q => 
                           REGISTERS_2_10_port, QN => n10595);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n11990, CK => n872, Q => 
                           REGISTERS_3_10_port, QN => n10627);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n12022, CK => n872, Q => 
                           REGISTERS_4_10_port, QN => n10659);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n12054, CK => n872, Q => 
                           REGISTERS_5_10_port, QN => n10691);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n12086, CK => n871, Q => 
                           REGISTERS_6_10_port, QN => n10723);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n12118, CK => n871, Q => 
                           REGISTERS_7_10_port, QN => n10755);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n12150, CK => n871, Q => 
                           REGISTERS_8_10_port, QN => n10787);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n12182, CK => n871, Q => 
                           REGISTERS_9_10_port, QN => n10819);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n12214_port, CK => n871, Q 
                           => REGISTERS_10_10_port, QN => n10851);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n12246_port, CK => n871, Q 
                           => REGISTERS_11_10_port, QN => n10883);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n12278_port, CK => n871, Q 
                           => REGISTERS_12_10_port, QN => n10915);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n12310, CK => n871, Q => 
                           REGISTERS_13_10_port, QN => n10947);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n12342, CK => n871, Q => 
                           REGISTERS_14_10_port, QN => n10979);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n12374, CK => n871, Q => 
                           REGISTERS_15_10_port, QN => n11011);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n12406, CK => n871, Q => 
                           REGISTERS_16_10_port, QN => n11043);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n12438, CK => n870, Q => 
                           REGISTERS_17_10_port, QN => n11075);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n12470, CK => n870, Q => 
                           REGISTERS_18_10_port, QN => n11107);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n12502, CK => n870, Q => 
                           REGISTERS_19_10_port, QN => n11139);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n12534, CK => n870, Q => 
                           REGISTERS_20_10_port, QN => n11171);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n12566, CK => n870, Q => 
                           REGISTERS_21_10_port, QN => n11203);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n12598, CK => n870, Q => 
                           REGISTERS_22_10_port, QN => n11235);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n12630, CK => n870, Q => 
                           REGISTERS_23_10_port, QN => n11267);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n12662, CK => n870, Q => 
                           REGISTERS_24_10_port, QN => n11299);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n12694, CK => n870, Q => 
                           REGISTERS_25_10_port, QN => n11331);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n12726, CK => n870, Q => 
                           REGISTERS_26_10_port, QN => n11363);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n12758, CK => n870, Q => 
                           REGISTERS_27_10_port, QN => n11395);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n12790, CK => n869, Q => 
                           REGISTERS_28_10_port, QN => n11427);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n12822, CK => n869, Q => 
                           REGISTERS_29_10_port, QN => n11459);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n12854, CK => n869, Q => 
                           REGISTERS_30_10_port, QN => n11491);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n12886, CK => n869, Q => 
                           REGISTERS_31_10_port, QN => n11523);
   REGISTERS_reg_32_10_inst : DFF_X1 port map( D => n12918, CK => n869, Q => 
                           REGISTERS_32_10_port, QN => n11555);
   REGISTERS_reg_33_10_inst : DFF_X1 port map( D => n12950, CK => n869, Q => 
                           REGISTERS_33_10_port, QN => n11587);
   REGISTERS_reg_34_10_inst : DFF_X1 port map( D => n12982, CK => n869, Q => 
                           REGISTERS_34_10_port, QN => n11619);
   REGISTERS_reg_35_10_inst : DFF_X1 port map( D => n13014, CK => n869, Q => 
                           REGISTERS_35_10_port, QN => n11651);
   REGISTERS_reg_36_10_inst : DFF_X1 port map( D => n13046, CK => n872, Q => 
                           REGISTERS_36_10_port, QN => n11683);
   REGISTERS_reg_38_9_inst : DFF_X1 port map( D => n13111, CK => n952, Q => 
                           REGISTERS_38_9_port, QN => n11748);
   REGISTERS_reg_39_9_inst : DFF_X1 port map( D => n13143, CK => n952, Q => 
                           REGISTERS_39_9_port, QN => n11780);
   REGISTERS_reg_37_9_inst : DFF_X1 port map( D => n13079, CK => n952, Q => 
                           REGISTERS_37_9_port, QN => n11716);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n11895, CK => n952, Q => 
                           REGISTERS_0_9_port, QN => n10514);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n11927, CK => n952, Q => 
                           REGISTERS_1_9_port, QN => n10564);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n11959, CK => n952, Q => 
                           REGISTERS_2_9_port, QN => n10596);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n11991, CK => n952, Q => 
                           REGISTERS_3_9_port, QN => n10628);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n12023, CK => n952, Q => 
                           REGISTERS_4_9_port, QN => n10660);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n12055, CK => n952, Q => 
                           REGISTERS_5_9_port, QN => n10692);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n12087, CK => n952, Q => 
                           REGISTERS_6_9_port, QN => n10724);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n12119, CK => n952, Q => 
                           REGISTERS_7_9_port, QN => n10756);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n12151, CK => n951, Q => 
                           REGISTERS_8_9_port, QN => n10788);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n12183, CK => n951, Q => 
                           REGISTERS_9_9_port, QN => n10820);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n12215_port, CK => n951, Q 
                           => REGISTERS_10_9_port, QN => n10852);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n12247_port, CK => n951, Q 
                           => REGISTERS_11_9_port, QN => n10884);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n12279_port, CK => n951, Q 
                           => REGISTERS_12_9_port, QN => n10916);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n12311, CK => n951, Q => 
                           REGISTERS_13_9_port, QN => n10948);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n12343, CK => n951, Q => 
                           REGISTERS_14_9_port, QN => n10980);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n12375, CK => n951, Q => 
                           REGISTERS_15_9_port, QN => n11012);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n12407, CK => n951, Q => 
                           REGISTERS_16_9_port, QN => n11044);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n12439, CK => n951, Q => 
                           REGISTERS_17_9_port, QN => n11076);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n12471, CK => n951, Q => 
                           REGISTERS_18_9_port, QN => n11108);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n12503, CK => n950, Q => 
                           REGISTERS_19_9_port, QN => n11140);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n12535, CK => n950, Q => 
                           REGISTERS_20_9_port, QN => n11172);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n12567, CK => n950, Q => 
                           REGISTERS_21_9_port, QN => n11204);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n12599, CK => n950, Q => 
                           REGISTERS_22_9_port, QN => n11236);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n12631, CK => n950, Q => 
                           REGISTERS_23_9_port, QN => n11268);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n12663, CK => n950, Q => 
                           REGISTERS_24_9_port, QN => n11300);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n12695, CK => n950, Q => 
                           REGISTERS_25_9_port, QN => n11332);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n12727, CK => n950, Q => 
                           REGISTERS_26_9_port, QN => n11364);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n12759, CK => n950, Q => 
                           REGISTERS_27_9_port, QN => n11396);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n12791, CK => n950, Q => 
                           REGISTERS_28_9_port, QN => n11428);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n12823, CK => n950, Q => 
                           REGISTERS_29_9_port, QN => n11460);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n12855, CK => n949, Q => 
                           REGISTERS_30_9_port, QN => n11492);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n12887, CK => n949, Q => 
                           REGISTERS_31_9_port, QN => n11524);
   REGISTERS_reg_32_9_inst : DFF_X1 port map( D => n12919, CK => n949, Q => 
                           REGISTERS_32_9_port, QN => n11556);
   REGISTERS_reg_33_9_inst : DFF_X1 port map( D => n12951, CK => n949, Q => 
                           REGISTERS_33_9_port, QN => n11588);
   REGISTERS_reg_34_9_inst : DFF_X1 port map( D => n12983, CK => n949, Q => 
                           REGISTERS_34_9_port, QN => n11620);
   REGISTERS_reg_35_9_inst : DFF_X1 port map( D => n13015, CK => n949, Q => 
                           REGISTERS_35_9_port, QN => n11652);
   REGISTERS_reg_36_9_inst : DFF_X1 port map( D => n13047, CK => n953, Q => 
                           REGISTERS_36_9_port, QN => n11684);
   REGISTERS_reg_38_8_inst : DFF_X1 port map( D => n13112, CK => n887, Q => 
                           REGISTERS_38_8_port, QN => n11749);
   REGISTERS_reg_39_8_inst : DFF_X1 port map( D => n13144, CK => n888, Q => 
                           REGISTERS_39_8_port, QN => n11781);
   REGISTERS_reg_37_8_inst : DFF_X1 port map( D => n13080, CK => n887, Q => 
                           REGISTERS_37_8_port, QN => n11717);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n11896, CK => n887, Q => 
                           REGISTERS_0_8_port, QN => n10517);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n11928, CK => n887, Q => 
                           REGISTERS_1_8_port, QN => n10565);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n11960, CK => n887, Q => 
                           REGISTERS_2_8_port, QN => n10597);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n11992, CK => n887, Q => 
                           REGISTERS_3_8_port, QN => n10629);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n12024, CK => n887, Q => 
                           REGISTERS_4_8_port, QN => n10661);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n12056, CK => n887, Q => 
                           REGISTERS_5_8_port, QN => n10693);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n12088, CK => n887, Q => 
                           REGISTERS_6_8_port, QN => n10725);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n12120, CK => n887, Q => 
                           REGISTERS_7_8_port, QN => n10757);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n12152, CK => n887, Q => 
                           REGISTERS_8_8_port, QN => n10789);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n12184, CK => n886, Q => 
                           REGISTERS_9_8_port, QN => n10821);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n12216_port, CK => n886, Q 
                           => REGISTERS_10_8_port, QN => n10853);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n12248_port, CK => n886, Q 
                           => REGISTERS_11_8_port, QN => n10885);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n12280_port, CK => n886, Q 
                           => REGISTERS_12_8_port, QN => n10917);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n12312, CK => n886, Q => 
                           REGISTERS_13_8_port, QN => n10949);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n12344, CK => n886, Q => 
                           REGISTERS_14_8_port, QN => n10981);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n12376, CK => n886, Q => 
                           REGISTERS_15_8_port, QN => n11013);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n12408, CK => n886, Q => 
                           REGISTERS_16_8_port, QN => n11045);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n12440, CK => n886, Q => 
                           REGISTERS_17_8_port, QN => n11077);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n12472, CK => n886, Q => 
                           REGISTERS_18_8_port, QN => n11109);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n12504, CK => n886, Q => 
                           REGISTERS_19_8_port, QN => n11141);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n12536, CK => n885, Q => 
                           REGISTERS_20_8_port, QN => n11173);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n12568, CK => n885, Q => 
                           REGISTERS_21_8_port, QN => n11205);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n12600, CK => n885, Q => 
                           REGISTERS_22_8_port, QN => n11237);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n12632, CK => n885, Q => 
                           REGISTERS_23_8_port, QN => n11269);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n12664, CK => n885, Q => 
                           REGISTERS_24_8_port, QN => n11301);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n12696, CK => n885, Q => 
                           REGISTERS_25_8_port, QN => n11333);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n12728, CK => n885, Q => 
                           REGISTERS_26_8_port, QN => n11365);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n12760, CK => n885, Q => 
                           REGISTERS_27_8_port, QN => n11397);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n12792, CK => n885, Q => 
                           REGISTERS_28_8_port, QN => n11429);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n12824, CK => n885, Q => 
                           REGISTERS_29_8_port, QN => n11461);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n12856, CK => n885, Q => 
                           REGISTERS_30_8_port, QN => n11493);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n12888, CK => n884, Q => 
                           REGISTERS_31_8_port, QN => n11525);
   REGISTERS_reg_32_8_inst : DFF_X1 port map( D => n12920, CK => n884, Q => 
                           REGISTERS_32_8_port, QN => n11557);
   REGISTERS_reg_33_8_inst : DFF_X1 port map( D => n12952, CK => n884, Q => 
                           REGISTERS_33_8_port, QN => n11589);
   REGISTERS_reg_34_8_inst : DFF_X1 port map( D => n12984, CK => n884, Q => 
                           REGISTERS_34_8_port, QN => n11621);
   REGISTERS_reg_35_8_inst : DFF_X1 port map( D => n13016, CK => n884, Q => 
                           REGISTERS_35_8_port, QN => n11653);
   REGISTERS_reg_36_8_inst : DFF_X1 port map( D => n13048, CK => n888, Q => 
                           REGISTERS_36_8_port, QN => n11685);
   REGISTERS_reg_38_7_inst : DFF_X1 port map( D => n13113, CK => n868, Q => 
                           REGISTERS_38_7_port, QN => n11750);
   REGISTERS_reg_39_7_inst : DFF_X1 port map( D => n13145, CK => n868, Q => 
                           REGISTERS_39_7_port, QN => n11782);
   REGISTERS_reg_37_7_inst : DFF_X1 port map( D => n13081, CK => n868, Q => 
                           REGISTERS_37_7_port, QN => n11718);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n11897, CK => n868, Q => 
                           REGISTERS_0_7_port, QN => n10520);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n11929, CK => n868, Q => 
                           REGISTERS_1_7_port, QN => n10566);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n11961, CK => n868, Q => 
                           REGISTERS_2_7_port, QN => n10598);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n11993, CK => n868, Q => 
                           REGISTERS_3_7_port, QN => n10630);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n12025, CK => n868, Q => 
                           REGISTERS_4_7_port, QN => n10662);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n12057, CK => n868, Q => 
                           REGISTERS_5_7_port, QN => n10694);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n12089, CK => n868, Q => 
                           REGISTERS_6_7_port, QN => n10726);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n12121, CK => n868, Q => 
                           REGISTERS_7_7_port, QN => n10758);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n12153, CK => n867, Q => 
                           REGISTERS_8_7_port, QN => n10790);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n12185, CK => n867, Q => 
                           REGISTERS_9_7_port, QN => n10822);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n12217_port, CK => n867, Q 
                           => REGISTERS_10_7_port, QN => n10854);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n12249_port, CK => n867, Q 
                           => REGISTERS_11_7_port, QN => n10886);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n12281_port, CK => n867, Q 
                           => REGISTERS_12_7_port, QN => n10918);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n12313, CK => n867, Q => 
                           REGISTERS_13_7_port, QN => n10950);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n12345, CK => n867, Q => 
                           REGISTERS_14_7_port, QN => n10982);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n12377, CK => n867, Q => 
                           REGISTERS_15_7_port, QN => n11014);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n12409, CK => n867, Q => 
                           REGISTERS_16_7_port, QN => n11046);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n12441, CK => n867, Q => 
                           REGISTERS_17_7_port, QN => n11078);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n12473, CK => n867, Q => 
                           REGISTERS_18_7_port, QN => n11110);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n12505, CK => n866, Q => 
                           REGISTERS_19_7_port, QN => n11142);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n12537, CK => n866, Q => 
                           REGISTERS_20_7_port, QN => n11174);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n12569, CK => n866, Q => 
                           REGISTERS_21_7_port, QN => n11206);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n12601, CK => n866, Q => 
                           REGISTERS_22_7_port, QN => n11238);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n12633, CK => n866, Q => 
                           REGISTERS_23_7_port, QN => n11270);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n12665, CK => n866, Q => 
                           REGISTERS_24_7_port, QN => n11302);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n12697, CK => n866, Q => 
                           REGISTERS_25_7_port, QN => n11334);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n12729, CK => n866, Q => 
                           REGISTERS_26_7_port, QN => n11366);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n12761, CK => n866, Q => 
                           REGISTERS_27_7_port, QN => n11398);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n12793, CK => n866, Q => 
                           REGISTERS_28_7_port, QN => n11430);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n12825, CK => n866, Q => 
                           REGISTERS_29_7_port, QN => n11462);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n12857, CK => n865, Q => 
                           REGISTERS_30_7_port, QN => n11494);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n12889, CK => n865, Q => 
                           REGISTERS_31_7_port, QN => n11526);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n12921, CK => n865, Q => 
                           REGISTERS_32_7_port, QN => n11558);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n12953, CK => n865, Q => 
                           REGISTERS_33_7_port, QN => n11590);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n12985, CK => n865, Q => 
                           REGISTERS_34_7_port, QN => n11622);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n13017, CK => n865, Q => 
                           REGISTERS_35_7_port, QN => n11654);
   REGISTERS_reg_36_7_inst : DFF_X1 port map( D => n13049, CK => n869, Q => 
                           REGISTERS_36_7_port, QN => n11686);
   REGISTERS_reg_38_6_inst : DFF_X1 port map( D => n13114, CK => n865, Q => 
                           REGISTERS_38_6_port, QN => n11751);
   REGISTERS_reg_39_6_inst : DFF_X1 port map( D => n13146, CK => n865, Q => 
                           REGISTERS_39_6_port, QN => n11783);
   REGISTERS_reg_37_6_inst : DFF_X1 port map( D => n13082, CK => n864, Q => 
                           REGISTERS_37_6_port, QN => n11719);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n11898, CK => n864, Q => 
                           REGISTERS_0_6_port, QN => n10523);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n11930, CK => n864, Q => 
                           REGISTERS_1_6_port, QN => n10567);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n11962, CK => n864, Q => 
                           REGISTERS_2_6_port, QN => n10599);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n11994, CK => n864, Q => 
                           REGISTERS_3_6_port, QN => n10631);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n12026, CK => n864, Q => 
                           REGISTERS_4_6_port, QN => n10663);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n12058, CK => n864, Q => 
                           REGISTERS_5_6_port, QN => n10695);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n12090, CK => n864, Q => 
                           REGISTERS_6_6_port, QN => n10727);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n12122, CK => n864, Q => 
                           REGISTERS_7_6_port, QN => n10759);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n12154, CK => n864, Q => 
                           REGISTERS_8_6_port, QN => n10791);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n12186, CK => n864, Q => 
                           REGISTERS_9_6_port, QN => n10823);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n12218_port, CK => n863, Q 
                           => REGISTERS_10_6_port, QN => n10855);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n12250_port, CK => n863, Q 
                           => REGISTERS_11_6_port, QN => n10887);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n12282_port, CK => n863, Q 
                           => REGISTERS_12_6_port, QN => n10919);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n12314, CK => n863, Q => 
                           REGISTERS_13_6_port, QN => n10951);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n12346, CK => n863, Q => 
                           REGISTERS_14_6_port, QN => n10983);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n12378, CK => n863, Q => 
                           REGISTERS_15_6_port, QN => n11015);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n12410, CK => n863, Q => 
                           REGISTERS_16_6_port, QN => n11047);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n12442, CK => n863, Q => 
                           REGISTERS_17_6_port, QN => n11079);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n12474, CK => n863, Q => 
                           REGISTERS_18_6_port, QN => n11111);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n12506, CK => n863, Q => 
                           REGISTERS_19_6_port, QN => n11143);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n12538, CK => n863, Q => 
                           REGISTERS_20_6_port, QN => n11175);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n12570, CK => n862, Q => 
                           REGISTERS_21_6_port, QN => n11207);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n12602, CK => n862, Q => 
                           REGISTERS_22_6_port, QN => n11239);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n12634, CK => n862, Q => 
                           REGISTERS_23_6_port, QN => n11271);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n12666, CK => n862, Q => 
                           REGISTERS_24_6_port, QN => n11303);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n12698, CK => n862, Q => 
                           REGISTERS_25_6_port, QN => n11335);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n12730, CK => n862, Q => 
                           REGISTERS_26_6_port, QN => n11367);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n12762, CK => n862, Q => 
                           REGISTERS_27_6_port, QN => n11399);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n12794, CK => n862, Q => 
                           REGISTERS_28_6_port, QN => n11431);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n12826, CK => n862, Q => 
                           REGISTERS_29_6_port, QN => n11463);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n12858, CK => n862, Q => 
                           REGISTERS_30_6_port, QN => n11495);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n12890, CK => n862, Q => 
                           REGISTERS_31_6_port, QN => n11527);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n12922, CK => n861, Q => 
                           REGISTERS_32_6_port, QN => n11559);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n12954, CK => n861, Q => 
                           REGISTERS_33_6_port, QN => n11591);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n12986, CK => n861, Q => 
                           REGISTERS_34_6_port, QN => n11623);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n13018, CK => n861, Q => 
                           REGISTERS_35_6_port, QN => n11655);
   REGISTERS_reg_36_6_inst : DFF_X1 port map( D => n13050, CK => n865, Q => 
                           REGISTERS_36_6_port, QN => n11687);
   REGISTERS_reg_38_5_inst : DFF_X1 port map( D => n13115, CK => n891, Q => 
                           REGISTERS_38_5_port, QN => n11752);
   REGISTERS_reg_39_5_inst : DFF_X1 port map( D => n13147, CK => n891, Q => 
                           REGISTERS_39_5_port, QN => n11784);
   REGISTERS_reg_37_5_inst : DFF_X1 port map( D => n13083, CK => n891, Q => 
                           REGISTERS_37_5_port, QN => n11720);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n11899, CK => n891, Q => 
                           REGISTERS_0_5_port, QN => n10526);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n11931, CK => n891, Q => 
                           REGISTERS_1_5_port, QN => n10568);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n11963, CK => n891, Q => 
                           REGISTERS_2_5_port, QN => n10600);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n11995, CK => n891, Q => 
                           REGISTERS_3_5_port, QN => n10632);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n12027, CK => n891, Q => 
                           REGISTERS_4_5_port, QN => n10664);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n12059, CK => n891, Q => 
                           REGISTERS_5_5_port, QN => n10696);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n12091, CK => n891, Q => 
                           REGISTERS_6_5_port, QN => n10728);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n12123, CK => n890, Q => 
                           REGISTERS_7_5_port, QN => n10760);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n12155, CK => n890, Q => 
                           REGISTERS_8_5_port, QN => n10792);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n12187, CK => n890, Q => 
                           REGISTERS_9_5_port, QN => n10824);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n12219_port, CK => n890, Q 
                           => REGISTERS_10_5_port, QN => n10856);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n12251_port, CK => n890, Q 
                           => REGISTERS_11_5_port, QN => n10888);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n12283_port, CK => n890, Q 
                           => REGISTERS_12_5_port, QN => n10920);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n12315, CK => n890, Q => 
                           REGISTERS_13_5_port, QN => n10952);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n12347, CK => n890, Q => 
                           REGISTERS_14_5_port, QN => n10984);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n12379, CK => n890, Q => 
                           REGISTERS_15_5_port, QN => n11016);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n12411, CK => n890, Q => 
                           REGISTERS_16_5_port, QN => n11048);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n12443, CK => n890, Q => 
                           REGISTERS_17_5_port, QN => n11080);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n12475, CK => n889, Q => 
                           REGISTERS_18_5_port, QN => n11112);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n12507, CK => n889, Q => 
                           REGISTERS_19_5_port, QN => n11144);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n12539, CK => n889, Q => 
                           REGISTERS_20_5_port, QN => n11176);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n12571, CK => n889, Q => 
                           REGISTERS_21_5_port, QN => n11208);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n12603, CK => n889, Q => 
                           REGISTERS_22_5_port, QN => n11240);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n12635, CK => n889, Q => 
                           REGISTERS_23_5_port, QN => n11272);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n12667, CK => n889, Q => 
                           REGISTERS_24_5_port, QN => n11304);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n12699, CK => n889, Q => 
                           REGISTERS_25_5_port, QN => n11336);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n12731, CK => n889, Q => 
                           REGISTERS_26_5_port, QN => n11368);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n12763, CK => n889, Q => 
                           REGISTERS_27_5_port, QN => n11400);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n12795, CK => n889, Q => 
                           REGISTERS_28_5_port, QN => n11432);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n12827, CK => n888, Q => 
                           REGISTERS_29_5_port, QN => n11464);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n12859, CK => n888, Q => 
                           REGISTERS_30_5_port, QN => n11496);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n12891, CK => n888, Q => 
                           REGISTERS_31_5_port, QN => n11528);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n12923, CK => n888, Q => 
                           REGISTERS_32_5_port, QN => n11560);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n12955, CK => n888, Q => 
                           REGISTERS_33_5_port, QN => n11592);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n12987, CK => n888, Q => 
                           REGISTERS_34_5_port, QN => n11624);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n13019, CK => n888, Q => 
                           REGISTERS_35_5_port, QN => n11656);
   REGISTERS_reg_36_5_inst : DFF_X1 port map( D => n13051, CK => n891, Q => 
                           REGISTERS_36_5_port, QN => n11688);
   REGISTERS_reg_38_4_inst : DFF_X1 port map( D => n13116, CK => n968, Q => 
                           REGISTERS_38_4_port, QN => n11753);
   REGISTERS_reg_39_4_inst : DFF_X1 port map( D => n13148, CK => n968, Q => 
                           REGISTERS_39_4_port, QN => n11785);
   REGISTERS_reg_37_4_inst : DFF_X1 port map( D => n13084, CK => n968, Q => 
                           REGISTERS_37_4_port, QN => n11721);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n11900, CK => n967, Q => 
                           REGISTERS_0_4_port, QN => n10529);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n11932, CK => n967, Q => 
                           REGISTERS_1_4_port, QN => n10569);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n11964, CK => n967, Q => 
                           REGISTERS_2_4_port, QN => n10601);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n11996, CK => n967, Q => 
                           REGISTERS_3_4_port, QN => n10633);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n12028, CK => n967, Q => 
                           REGISTERS_4_4_port, QN => n10665);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n12060, CK => n967, Q => 
                           REGISTERS_5_4_port, QN => n10697);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n12092, CK => n967, Q => 
                           REGISTERS_6_4_port, QN => n10729);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n12124, CK => n967, Q => 
                           REGISTERS_7_4_port, QN => n10761);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n12156, CK => n967, Q => 
                           REGISTERS_8_4_port, QN => n10793);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n12188, CK => n967, Q => 
                           REGISTERS_9_4_port, QN => n10825);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n12220_port, CK => n967, Q 
                           => REGISTERS_10_4_port, QN => n10857);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n12252_port, CK => n966, Q 
                           => REGISTERS_11_4_port, QN => n10889);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n12284_port, CK => n966, Q 
                           => REGISTERS_12_4_port, QN => n10921);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n12316, CK => n966, Q => 
                           REGISTERS_13_4_port, QN => n10953);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n12348, CK => n966, Q => 
                           REGISTERS_14_4_port, QN => n10985);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n12380, CK => n966, Q => 
                           REGISTERS_15_4_port, QN => n11017);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n12412, CK => n966, Q => 
                           REGISTERS_16_4_port, QN => n11049);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n12444, CK => n966, Q => 
                           REGISTERS_17_4_port, QN => n11081);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n12476, CK => n966, Q => 
                           REGISTERS_18_4_port, QN => n11113);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n12508, CK => n966, Q => 
                           REGISTERS_19_4_port, QN => n11145);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n12540, CK => n966, Q => 
                           REGISTERS_20_4_port, QN => n11177);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n12572, CK => n966, Q => 
                           REGISTERS_21_4_port, QN => n11209);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n12604, CK => n965, Q => 
                           REGISTERS_22_4_port, QN => n11241);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n12636, CK => n965, Q => 
                           REGISTERS_23_4_port, QN => n11273);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n12668, CK => n965, Q => 
                           REGISTERS_24_4_port, QN => n11305);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n12700, CK => n965, Q => 
                           REGISTERS_25_4_port, QN => n11337);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n12732, CK => n965, Q => 
                           REGISTERS_26_4_port, QN => n11369);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n12764, CK => n965, Q => 
                           REGISTERS_27_4_port, QN => n11401);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n12796, CK => n965, Q => 
                           REGISTERS_28_4_port, QN => n11433);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n12828, CK => n965, Q => 
                           REGISTERS_29_4_port, QN => n11465);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n12860, CK => n965, Q => 
                           REGISTERS_30_4_port, QN => n11497);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n12892, CK => n965, Q => 
                           REGISTERS_31_4_port, QN => n11529);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n12924, CK => n965, Q => 
                           REGISTERS_32_4_port, QN => n11561);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n12956, CK => n964, Q => 
                           REGISTERS_33_4_port, QN => n11593);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n12988, CK => n964, Q => 
                           REGISTERS_34_4_port, QN => n11625);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n13020, CK => n964, Q => 
                           REGISTERS_35_4_port, QN => n11657);
   REGISTERS_reg_36_4_inst : DFF_X1 port map( D => n13052, CK => n968, Q => 
                           REGISTERS_36_4_port, QN => n11689);
   REGISTERS_reg_38_3_inst : DFF_X1 port map( D => n13117, CK => n861, Q => 
                           REGISTERS_38_3_port, QN => n11754);
   REGISTERS_reg_39_3_inst : DFF_X1 port map( D => n13149, CK => n861, Q => 
                           REGISTERS_39_3_port, QN => n11786);
   REGISTERS_reg_37_3_inst : DFF_X1 port map( D => n13085, CK => n861, Q => 
                           REGISTERS_37_3_port, QN => n11722);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n11901, CK => n861, Q => 
                           REGISTERS_0_3_port, QN => n10532);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n11933, CK => n860, Q => 
                           REGISTERS_1_3_port, QN => n10570);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n11965, CK => n860, Q => 
                           REGISTERS_2_3_port, QN => n10602);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n11997, CK => n860, Q => 
                           REGISTERS_3_3_port, QN => n10634);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n12029, CK => n860, Q => 
                           REGISTERS_4_3_port, QN => n10666);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n12061, CK => n860, Q => 
                           REGISTERS_5_3_port, QN => n10698);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n12093, CK => n860, Q => 
                           REGISTERS_6_3_port, QN => n10730);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n12125, CK => n860, Q => 
                           REGISTERS_7_3_port, QN => n10762);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n12157, CK => n860, Q => 
                           REGISTERS_8_3_port, QN => n10794);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n12189, CK => n860, Q => 
                           REGISTERS_9_3_port, QN => n10826);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n12221_port, CK => n860, Q 
                           => REGISTERS_10_3_port, QN => n10858);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n12253_port, CK => n860, Q 
                           => REGISTERS_11_3_port, QN => n10890);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n12285_port, CK => n859, Q 
                           => REGISTERS_12_3_port, QN => n10922);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n12317, CK => n859, Q => 
                           REGISTERS_13_3_port, QN => n10954);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n12349, CK => n859, Q => 
                           REGISTERS_14_3_port, QN => n10986);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n12381, CK => n859, Q => 
                           REGISTERS_15_3_port, QN => n11018);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n12413, CK => n859, Q => 
                           REGISTERS_16_3_port, QN => n11050);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n12445, CK => n859, Q => 
                           REGISTERS_17_3_port, QN => n11082);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n12477, CK => n859, Q => 
                           REGISTERS_18_3_port, QN => n11114);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n12509, CK => n859, Q => 
                           REGISTERS_19_3_port, QN => n11146);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n12541, CK => n859, Q => 
                           REGISTERS_20_3_port, QN => n11178);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n12573, CK => n859, Q => 
                           REGISTERS_21_3_port, QN => n11210);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n12605, CK => n859, Q => 
                           REGISTERS_22_3_port, QN => n11242);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n12637, CK => n858, Q => 
                           REGISTERS_23_3_port, QN => n11274);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n12669, CK => n858, Q => 
                           REGISTERS_24_3_port, QN => n11306);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n12701, CK => n858, Q => 
                           REGISTERS_25_3_port, QN => n11338);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n12733, CK => n858, Q => 
                           REGISTERS_26_3_port, QN => n11370);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n12765, CK => n858, Q => 
                           REGISTERS_27_3_port, QN => n11402);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n12797, CK => n858, Q => 
                           REGISTERS_28_3_port, QN => n11434);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n12829, CK => n858, Q => 
                           REGISTERS_29_3_port, QN => n11466);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n12861, CK => n858, Q => 
                           REGISTERS_30_3_port, QN => n11498);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n12893, CK => n858, Q => 
                           REGISTERS_31_3_port, QN => n11530);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n12925, CK => n858, Q => 
                           REGISTERS_32_3_port, QN => n11562);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n12957, CK => n858, Q => 
                           REGISTERS_33_3_port, QN => n11594);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n12989, CK => n857, Q => 
                           REGISTERS_34_3_port, QN => n11626);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n13021, CK => n857, Q => 
                           REGISTERS_35_3_port, QN => n11658);
   REGISTERS_reg_36_3_inst : DFF_X1 port map( D => n13053, CK => n861, Q => 
                           REGISTERS_36_3_port, QN => n11690);
   REGISTERS_reg_38_2_inst : DFF_X1 port map( D => n13118, CK => n857, Q => 
                           REGISTERS_38_2_port, QN => n11755);
   REGISTERS_reg_39_2_inst : DFF_X1 port map( D => n13150, CK => n857, Q => 
                           REGISTERS_39_2_port, QN => n11787);
   REGISTERS_reg_37_2_inst : DFF_X1 port map( D => n13086, CK => n857, Q => 
                           REGISTERS_37_2_port, QN => n11723);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n11902, CK => n857, Q => 
                           REGISTERS_0_2_port, QN => n10535);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n11934, CK => n857, Q => 
                           REGISTERS_1_2_port, QN => n10571);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n11966, CK => n857, Q => 
                           REGISTERS_2_2_port, QN => n10603);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n11998, CK => n856, Q => 
                           REGISTERS_3_2_port, QN => n10635);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n12030, CK => n856, Q => 
                           REGISTERS_4_2_port, QN => n10667);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n12062, CK => n856, Q => 
                           REGISTERS_5_2_port, QN => n10699);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n12094, CK => n856, Q => 
                           REGISTERS_6_2_port, QN => n10731);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n12126, CK => n856, Q => 
                           REGISTERS_7_2_port, QN => n10763);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n12158, CK => n856, Q => 
                           REGISTERS_8_2_port, QN => n10795);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n12190, CK => n856, Q => 
                           REGISTERS_9_2_port, QN => n10827);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n12222_port, CK => n856, Q 
                           => REGISTERS_10_2_port, QN => n10859);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n12254_port, CK => n856, Q 
                           => REGISTERS_11_2_port, QN => n10891);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n12286_port, CK => n856, Q 
                           => REGISTERS_12_2_port, QN => n10923);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n12318, CK => n856, Q => 
                           REGISTERS_13_2_port, QN => n10955);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n12350, CK => n855, Q => 
                           REGISTERS_14_2_port, QN => n10987);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n12382, CK => n855, Q => 
                           REGISTERS_15_2_port, QN => n11019);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n12414, CK => n855, Q => 
                           REGISTERS_16_2_port, QN => n11051);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n12446, CK => n855, Q => 
                           REGISTERS_17_2_port, QN => n11083);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n12478, CK => n855, Q => 
                           REGISTERS_18_2_port, QN => n11115);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n12510, CK => n855, Q => 
                           REGISTERS_19_2_port, QN => n11147);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n12542, CK => n855, Q => 
                           REGISTERS_20_2_port, QN => n11179);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n12574, CK => n855, Q => 
                           REGISTERS_21_2_port, QN => n11211);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n12606, CK => n855, Q => 
                           REGISTERS_22_2_port, QN => n11243);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n12638, CK => n855, Q => 
                           REGISTERS_23_2_port, QN => n11275);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n12670, CK => n855, Q => 
                           REGISTERS_24_2_port, QN => n11307);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n12702, CK => n854, Q => 
                           REGISTERS_25_2_port, QN => n11339);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n12734, CK => n854, Q => 
                           REGISTERS_26_2_port, QN => n11371);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n12766, CK => n854, Q => 
                           REGISTERS_27_2_port, QN => n11403);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n12798, CK => n854, Q => 
                           REGISTERS_28_2_port, QN => n11435);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n12830, CK => n854, Q => 
                           REGISTERS_29_2_port, QN => n11467);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n12862, CK => n854, Q => 
                           REGISTERS_30_2_port, QN => n11499);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n12894, CK => n854, Q => 
                           REGISTERS_31_2_port, QN => n11531);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n12926, CK => n854, Q => 
                           REGISTERS_32_2_port, QN => n11563);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n12958, CK => n854, Q => 
                           REGISTERS_33_2_port, QN => n11595);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n12990, CK => n854, Q => 
                           REGISTERS_34_2_port, QN => n11627);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n13022, CK => n854, Q => 
                           REGISTERS_35_2_port, QN => n11659);
   REGISTERS_reg_36_2_inst : DFF_X1 port map( D => n13054, CK => n857, Q => 
                           REGISTERS_36_2_port, QN => n11691);
   REGISTERS_reg_38_1_inst : DFF_X1 port map( D => n13119, CK => n853, Q => 
                           REGISTERS_38_1_port, QN => n11756);
   REGISTERS_reg_39_1_inst : DFF_X1 port map( D => n13151, CK => n853, Q => 
                           REGISTERS_39_1_port, QN => n11788);
   REGISTERS_reg_37_1_inst : DFF_X1 port map( D => n13087, CK => n853, Q => 
                           REGISTERS_37_1_port, QN => n11724);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n11903, CK => n853, Q => 
                           REGISTERS_0_1_port, QN => n10538);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n11935, CK => n853, Q => 
                           REGISTERS_1_1_port, QN => n10572);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n11967, CK => n853, Q => 
                           REGISTERS_2_1_port, QN => n10604);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n11999, CK => n853, Q => 
                           REGISTERS_3_1_port, QN => n10636);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n12031, CK => n853, Q => 
                           REGISTERS_4_1_port, QN => n10668);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n12063, CK => n852, Q => 
                           REGISTERS_5_1_port, QN => n10700);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n12095, CK => n852, Q => 
                           REGISTERS_6_1_port, QN => n10732);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n12127, CK => n852, Q => 
                           REGISTERS_7_1_port, QN => n10764);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n12159, CK => n852, Q => 
                           REGISTERS_8_1_port, QN => n10796);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n12191, CK => n852, Q => 
                           REGISTERS_9_1_port, QN => n10828);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n12223_port, CK => n852, Q 
                           => REGISTERS_10_1_port, QN => n10860);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n12255_port, CK => n852, Q 
                           => REGISTERS_11_1_port, QN => n10892);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n12287_port, CK => n852, Q 
                           => REGISTERS_12_1_port, QN => n10924);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n12319, CK => n852, Q => 
                           REGISTERS_13_1_port, QN => n10956);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n12351, CK => n852, Q => 
                           REGISTERS_14_1_port, QN => n10988);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n12383, CK => n852, Q => 
                           REGISTERS_15_1_port, QN => n11020);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n12415, CK => n851, Q => 
                           REGISTERS_16_1_port, QN => n11052);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n12447, CK => n851, Q => 
                           REGISTERS_17_1_port, QN => n11084);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n12479, CK => n851, Q => 
                           REGISTERS_18_1_port, QN => n11116);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n12511, CK => n851, Q => 
                           REGISTERS_19_1_port, QN => n11148);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n12543, CK => n851, Q => 
                           REGISTERS_20_1_port, QN => n11180);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n12575, CK => n851, Q => 
                           REGISTERS_21_1_port, QN => n11212);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n12607, CK => n851, Q => 
                           REGISTERS_22_1_port, QN => n11244);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n12639, CK => n851, Q => 
                           REGISTERS_23_1_port, QN => n11276);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n12671, CK => n851, Q => 
                           REGISTERS_24_1_port, QN => n11308);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n12703, CK => n851, Q => 
                           REGISTERS_25_1_port, QN => n11340);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n12735, CK => n851, Q => 
                           REGISTERS_26_1_port, QN => n11372);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n12767, CK => n850, Q => 
                           REGISTERS_27_1_port, QN => n11404);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n12799, CK => n850, Q => 
                           REGISTERS_28_1_port, QN => n11436);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n12831, CK => n850, Q => 
                           REGISTERS_29_1_port, QN => n11468);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n12863, CK => n850, Q => 
                           REGISTERS_30_1_port, QN => n11500);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n12895, CK => n850, Q => 
                           REGISTERS_31_1_port, QN => n11532);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n12927, CK => n850, Q => 
                           REGISTERS_32_1_port, QN => n11564);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n12959, CK => n850, Q => 
                           REGISTERS_33_1_port, QN => n11596);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n12991, CK => n850, Q => 
                           REGISTERS_34_1_port, QN => n11628);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n13023, CK => n850, Q => 
                           REGISTERS_35_1_port, QN => n11660);
   REGISTERS_reg_36_1_inst : DFF_X1 port map( D => n13055, CK => n853, Q => 
                           REGISTERS_36_1_port, QN => n11692);
   REGISTERS_reg_38_0_inst : DFF_X1 port map( D => n13120, CK => n971, Q => 
                           REGISTERS_38_0_port, QN => n11757);
   REGISTERS_reg_39_0_inst : DFF_X1 port map( D => n13152, CK => n971, Q => 
                           REGISTERS_39_0_port, QN => n11789);
   REGISTERS_reg_37_0_inst : DFF_X1 port map( D => n13088, CK => n971, Q => 
                           REGISTERS_37_0_port, QN => n11725);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n11904, CK => n971, Q => 
                           REGISTERS_0_0_port, QN => n10541);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n11936, CK => n971, Q => 
                           REGISTERS_1_0_port, QN => n10573);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n11968, CK => n971, Q => 
                           REGISTERS_2_0_port, QN => n10605);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n12000, CK => n971, Q => 
                           REGISTERS_3_0_port, QN => n10637);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n12032, CK => n971, Q => 
                           REGISTERS_4_0_port, QN => n10669);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n12064, CK => n971, Q => 
                           REGISTERS_5_0_port, QN => n10701);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n12096, CK => n971, Q => 
                           REGISTERS_6_0_port, QN => n10733);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n12128, CK => n971, Q => 
                           REGISTERS_7_0_port, QN => n10765);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n12160, CK => n970, Q => 
                           REGISTERS_8_0_port, QN => n10797);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n12192, CK => n970, Q => 
                           REGISTERS_9_0_port, QN => n10829);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n12224_port, CK => n970, Q 
                           => REGISTERS_10_0_port, QN => n10861);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n12256_port, CK => n970, Q 
                           => REGISTERS_11_0_port, QN => n10893);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n12288_port, CK => n970, Q 
                           => REGISTERS_12_0_port, QN => n10925);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n12320, CK => n970, Q => 
                           REGISTERS_13_0_port, QN => n10957);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n12352, CK => n970, Q => 
                           REGISTERS_14_0_port, QN => n10989);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n12384, CK => n970, Q => 
                           REGISTERS_15_0_port, QN => n11021);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n12416, CK => n970, Q => 
                           REGISTERS_16_0_port, QN => n11053);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n12448, CK => n970, Q => 
                           REGISTERS_17_0_port, QN => n11085);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n12480, CK => n970, Q => 
                           REGISTERS_18_0_port, QN => n11117);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n12512, CK => n969, Q => 
                           REGISTERS_19_0_port, QN => n11149);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n12544, CK => n969, Q => 
                           REGISTERS_20_0_port, QN => n11181);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n12576, CK => n969, Q => 
                           REGISTERS_21_0_port, QN => n11213);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n12608, CK => n969, Q => 
                           REGISTERS_22_0_port, QN => n11245);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n12640, CK => n969, Q => 
                           REGISTERS_23_0_port, QN => n11277);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n12672, CK => n969, Q => 
                           REGISTERS_24_0_port, QN => n11309);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n12704, CK => n969, Q => 
                           REGISTERS_25_0_port, QN => n11341);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n12736, CK => n969, Q => 
                           REGISTERS_26_0_port, QN => n11373);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n12768, CK => n969, Q => 
                           REGISTERS_27_0_port, QN => n11405);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n12800, CK => n969, Q => 
                           REGISTERS_28_0_port, QN => n11437);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n12832, CK => n969, Q => 
                           REGISTERS_29_0_port, QN => n11469);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n12864, CK => n968, Q => 
                           REGISTERS_30_0_port, QN => n11501);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n12896, CK => n968, Q => 
                           REGISTERS_31_0_port, QN => n11533);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n12928, CK => n968, Q => 
                           REGISTERS_32_0_port, QN => n11565);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n12960, CK => n968, Q => 
                           REGISTERS_33_0_port, QN => n11597);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n12992, CK => n968, Q => 
                           REGISTERS_34_0_port, QN => n11629);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n13024, CK => n968, Q => 
                           REGISTERS_35_0_port, QN => n11661);
   REGISTERS_reg_36_0_inst : DFF_X1 port map( D => n13056, CK => n972, Q => 
                           REGISTERS_36_0_port, QN => n11693);
   REGISTERS_reg_39_31_inst : DFF_X1 port map( D => n13121, CK => n956, Q => 
                           REGISTERS_39_31_port, QN => n11758);
   REGISTERS_reg_38_31_inst : DFF_X1 port map( D => n13089, CK => n956, Q => 
                           REGISTERS_38_31_port, QN => n11726);
   REGISTERS_reg_36_31_inst : DFF_X1 port map( D => n13025, CK => n956, Q => 
                           REGISTERS_36_31_port, QN => n11662);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n11873, CK => n956, Q => 
                           REGISTERS_0_31_port, QN => n10448);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n11905, CK => n956, Q => 
                           REGISTERS_1_31_port, QN => n10542);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n11937, CK => n956, Q => 
                           REGISTERS_2_31_port, QN => n10574);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n11969, CK => n956, Q => 
                           REGISTERS_3_31_port, QN => n10606);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n12001, CK => n956, Q => 
                           REGISTERS_4_31_port, QN => n10638);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n12033, CK => n956, Q => 
                           REGISTERS_5_31_port, QN => n10670);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n12065, CK => n955, Q => 
                           REGISTERS_6_31_port, QN => n10702);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n12097, CK => n955, Q => 
                           REGISTERS_7_31_port, QN => n10734);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n12129, CK => n955, Q => 
                           REGISTERS_8_31_port, QN => n10766);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n12161, CK => n955, Q => 
                           REGISTERS_9_31_port, QN => n10798);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n12193, CK => n955, Q => 
                           REGISTERS_10_31_port, QN => n10830);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n12225_port, CK => n955, Q 
                           => REGISTERS_11_31_port, QN => n10862);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n12257_port, CK => n955, Q 
                           => REGISTERS_12_31_port, QN => n10894);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n12289_port, CK => n955, Q 
                           => REGISTERS_13_31_port, QN => n10926);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n12321, CK => n955, Q => 
                           REGISTERS_14_31_port, QN => n10958);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n12353, CK => n955, Q => 
                           REGISTERS_15_31_port, QN => n10990);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n12385, CK => n955, Q => 
                           REGISTERS_16_31_port, QN => n11022);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n12417, CK => n954, Q => 
                           REGISTERS_17_31_port, QN => n11054);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n12449, CK => n954, Q => 
                           REGISTERS_18_31_port, QN => n11086);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n12481, CK => n954, Q => 
                           REGISTERS_19_31_port, QN => n11118);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n12513, CK => n954, Q => 
                           REGISTERS_20_31_port, QN => n11150);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n12545, CK => n954, Q => 
                           REGISTERS_21_31_port, QN => n11182);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n12577, CK => n954, Q => 
                           REGISTERS_22_31_port, QN => n11214);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n12609, CK => n954, Q => 
                           REGISTERS_23_31_port, QN => n11246);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n12641, CK => n954, Q => 
                           REGISTERS_24_31_port, QN => n11278);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n12673, CK => n954, Q => 
                           REGISTERS_25_31_port, QN => n11310);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n12705, CK => n954, Q => 
                           REGISTERS_26_31_port, QN => n11342);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n12737, CK => n954, Q => 
                           REGISTERS_27_31_port, QN => n11374);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n12769, CK => n953, Q => 
                           REGISTERS_28_31_port, QN => n11406);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n12801, CK => n953, Q => 
                           REGISTERS_29_31_port, QN => n11438);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n12833, CK => n953, Q => 
                           REGISTERS_30_31_port, QN => n11470);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n12865, CK => n953, Q => 
                           REGISTERS_31_31_port, QN => n11502);
   REGISTERS_reg_32_31_inst : DFF_X1 port map( D => n12897, CK => n953, Q => 
                           REGISTERS_32_31_port, QN => n11534);
   REGISTERS_reg_33_31_inst : DFF_X1 port map( D => n12929, CK => n953, Q => 
                           REGISTERS_33_31_port, QN => n11566);
   REGISTERS_reg_34_31_inst : DFF_X1 port map( D => n12961, CK => n953, Q => 
                           REGISTERS_34_31_port, QN => n11598);
   REGISTERS_reg_35_31_inst : DFF_X1 port map( D => n12993, CK => n953, Q => 
                           REGISTERS_35_31_port, QN => n11630);
   REGISTERS_reg_37_31_inst : DFF_X1 port map( D => n13057, CK => n956, Q => 
                           REGISTERS_37_31_port, QN => n11694);
   MEM_OUT_reg_31_inst : DFF_X1 port map( D => n16456, CK => n981, Q => 
                           MEM_OUT_31_port, QN => n_1470);
   MEM_OUT_reg_30_inst : DFF_X1 port map( D => n16457, CK => n981, Q => 
                           MEM_OUT_30_port, QN => n_1471);
   MEM_OUT_reg_29_inst : DFF_X1 port map( D => n16458, CK => n980, Q => 
                           MEM_OUT_29_port, QN => n_1472);
   MEM_OUT_reg_28_inst : DFF_X1 port map( D => n16459, CK => n980, Q => 
                           MEM_OUT_28_port, QN => n_1473);
   MEM_OUT_reg_27_inst : DFF_X1 port map( D => n16460, CK => n980, Q => 
                           MEM_OUT_27_port, QN => n_1474);
   MEM_OUT_reg_26_inst : DFF_X1 port map( D => n16461, CK => n980, Q => 
                           MEM_OUT_26_port, QN => n_1475);
   MEM_OUT_reg_25_inst : DFF_X1 port map( D => n16462, CK => n980, Q => 
                           MEM_OUT_25_port, QN => n_1476);
   MEM_OUT_reg_24_inst : DFF_X1 port map( D => n16463, CK => n980, Q => 
                           MEM_OUT_24_port, QN => n_1477);
   MEM_OUT_reg_23_inst : DFF_X1 port map( D => n16464, CK => n980, Q => 
                           MEM_OUT_23_port, QN => n_1478);
   MEM_OUT_reg_22_inst : DFF_X1 port map( D => n16465, CK => n980, Q => 
                           MEM_OUT_22_port, QN => n_1479);
   MEM_OUT_reg_21_inst : DFF_X1 port map( D => n16466, CK => n980, Q => 
                           MEM_OUT_21_port, QN => n_1480);
   MEM_OUT_reg_20_inst : DFF_X1 port map( D => n16467, CK => n980, Q => 
                           MEM_OUT_20_port, QN => n_1481);
   MEM_OUT_reg_19_inst : DFF_X1 port map( D => n16468, CK => n980, Q => 
                           MEM_OUT_19_port, QN => n_1482);
   MEM_OUT_reg_18_inst : DFF_X1 port map( D => n16469, CK => n979, Q => 
                           MEM_OUT_18_port, QN => n_1483);
   MEM_OUT_reg_17_inst : DFF_X1 port map( D => n16470, CK => n979, Q => 
                           MEM_OUT_17_port, QN => n_1484);
   MEM_OUT_reg_16_inst : DFF_X1 port map( D => n16471, CK => n979, Q => 
                           MEM_OUT_16_port, QN => n_1485);
   MEM_OUT_reg_15_inst : DFF_X1 port map( D => n16472, CK => n979, Q => 
                           MEM_OUT_15_port, QN => n_1486);
   MEM_OUT_reg_14_inst : DFF_X1 port map( D => n16473, CK => n979, Q => 
                           MEM_OUT_14_port, QN => n_1487);
   MEM_OUT_reg_13_inst : DFF_X1 port map( D => n16474, CK => n979, Q => 
                           MEM_OUT_13_port, QN => n_1488);
   MEM_OUT_reg_12_inst : DFF_X1 port map( D => n16475, CK => n979, Q => 
                           MEM_OUT_12_port, QN => n_1489);
   MEM_OUT_reg_11_inst : DFF_X1 port map( D => n16476, CK => n979, Q => 
                           MEM_OUT_11_port, QN => n_1490);
   MEM_OUT_reg_10_inst : DFF_X1 port map( D => n16477, CK => n979, Q => 
                           MEM_OUT_10_port, QN => n_1491);
   MEM_OUT_reg_9_inst : DFF_X1 port map( D => n16478, CK => n979, Q => 
                           MEM_OUT_9_port, QN => n_1492);
   MEM_OUT_reg_8_inst : DFF_X1 port map( D => n16479, CK => n979, Q => 
                           MEM_OUT_8_port, QN => n_1493);
   MEM_OUT_reg_7_inst : DFF_X1 port map( D => n16480, CK => n978, Q => 
                           MEM_OUT_7_port, QN => n_1494);
   MEM_OUT_reg_6_inst : DFF_X1 port map( D => n16481, CK => n978, Q => 
                           MEM_OUT_6_port, QN => n_1495);
   MEM_OUT_reg_5_inst : DFF_X1 port map( D => n16482, CK => n978, Q => 
                           MEM_OUT_5_port, QN => n_1496);
   MEM_OUT_reg_4_inst : DFF_X1 port map( D => n16483, CK => n978, Q => 
                           MEM_OUT_4_port, QN => n_1497);
   MEM_OUT_reg_3_inst : DFF_X1 port map( D => n16484, CK => n978, Q => 
                           MEM_OUT_3_port, QN => n_1498);
   MEM_OUT_reg_2_inst : DFF_X1 port map( D => n16485, CK => n978, Q => 
                           MEM_OUT_2_port, QN => n_1499);
   MEM_OUT_reg_1_inst : DFF_X1 port map( D => n16486, CK => n978, Q => 
                           MEM_OUT_1_port, QN => n_1500);
   MEM_OUT_reg_0_inst : DFF_X1 port map( D => n16487, CK => n978, Q => 
                           MEM_OUT_0_port, QN => n_1501);
   FILL_reg : DFF_X1 port map( D => n11872, CK => n974, Q => FILL_port, QN => 
                           n_1502);
   n90 <= '1';
   n89 <= '0';
   SPILL <= '0';
   add_171 : window_rf_M4_N4_F4_NBIT32_DW01_add_0 port map( A(31) => 
                           SWP_31_port, A(30) => SWP_30_port, A(29) => 
                           SWP_29_port, A(28) => SWP_28_port, A(27) => 
                           SWP_27_port, A(26) => SWP_26_port, A(25) => 
                           SWP_25_port, A(24) => SWP_24_port, A(23) => 
                           SWP_23_port, A(22) => SWP_22_port, A(21) => 
                           SWP_21_port, A(20) => SWP_20_port, A(19) => 
                           SWP_19_port, A(18) => SWP_18_port, A(17) => 
                           SWP_17_port, A(16) => SWP_16_port, A(15) => 
                           SWP_15_port, A(14) => SWP_14_port, A(13) => 
                           SWP_13_port, A(12) => SWP_12_port, A(11) => 
                           SWP_11_port, A(10) => SWP_10_port, A(9) => 
                           SWP_9_port, A(8) => SWP_8_port, A(7) => SWP_7_port, 
                           A(6) => SWP_6_port, A(5) => n846, A(4) => n841, A(3)
                           => n302, A(2) => n301, A(1) => n840, A(0) => n804, 
                           B(31) => X_Logic0_port, B(30) => X_Logic0_port, 
                           B(29) => X_Logic0_port, B(28) => X_Logic0_port, 
                           B(27) => X_Logic0_port, B(26) => X_Logic0_port, 
                           B(25) => X_Logic0_port, B(24) => X_Logic0_port, 
                           B(23) => X_Logic0_port, B(22) => X_Logic0_port, 
                           B(21) => X_Logic0_port, B(20) => X_Logic0_port, 
                           B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
                           B(17) => X_Logic0_port, B(16) => X_Logic0_port, 
                           B(15) => X_Logic0_port, B(14) => X_Logic0_port, 
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic1_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, CI => n49, 
                           SUM(31) => N12268, SUM(30) => N12267, SUM(29) => 
                           N12266, SUM(28) => N12265, SUM(27) => N12264, 
                           SUM(26) => N12263, SUM(25) => N12262, SUM(24) => 
                           N12261, SUM(23) => N12260, SUM(22) => N12259, 
                           SUM(21) => N12258, SUM(20) => N12257, SUM(19) => 
                           N12256, SUM(18) => N12255, SUM(17) => N12254, 
                           SUM(16) => N12253, SUM(15) => N12252, SUM(14) => 
                           N12251, SUM(13) => N12250, SUM(12) => N12249, 
                           SUM(11) => N12248, SUM(10) => N12247, SUM(9) => 
                           N12246, SUM(8) => N12245, SUM(7) => N12244, SUM(6) 
                           => N12243, SUM(5) => N12242, SUM(4) => N12241, 
                           SUM(3) => N12240, SUM(2) => N12239, SUM(1) => N12238
                           , SUM(0) => N12237, CO => n_1503);
   add_65 : window_rf_M4_N4_F4_NBIT32_DW01_add_1 port map( A(5) => CWP_5_port, 
                           A(4) => CWP_4_port, A(3) => CWP_3_port, A(2) => 
                           CWP_2_port, A(1) => CWP_1_port, A(0) => CWP_0_port, 
                           B(5) => X_Logic0_port, B(4) => N3592, B(3) => N3591,
                           B(2) => N3590, B(1) => WR_ADD(1), B(0) => WR_ADD(0),
                           CI => n52, SUM(5) => N3598, SUM(4) => N3597, SUM(3) 
                           => N3596, SUM(2) => N3595, SUM(1) => N3594, SUM(0) 
                           => N3593, CO => n_1504);
   add_64 : window_rf_M4_N4_F4_NBIT32_DW01_add_2 port map( A(5) => CWP_5_port, 
                           A(4) => CWP_4_port, A(3) => CWP_3_port, A(2) => 
                           CWP_2_port, A(1) => CWP_1_port, A(0) => CWP_0_port, 
                           B(5) => X_Logic0_port, B(4) => N3579, B(3) => N3578,
                           B(2) => N3577, B(1) => RD2_ADD(1), B(0) => 
                           RD2_ADD(0), CI => n55, SUM(5) => N3585, SUM(4) => 
                           N3584, SUM(3) => N3583, SUM(2) => N3582, SUM(1) => 
                           N3581, SUM(0) => N3580, CO => n_1505);
   add_63 : window_rf_M4_N4_F4_NBIT32_DW01_add_3 port map( A(5) => CWP_5_port, 
                           A(4) => CWP_4_port, A(3) => CWP_3_port, A(2) => 
                           CWP_2_port, A(1) => CWP_1_port, A(0) => CWP_0_port, 
                           B(5) => X_Logic0_port, B(4) => N3566, B(3) => N3565,
                           B(2) => N3564, B(1) => RD1_ADD(1), B(0) => 
                           RD1_ADD(0), CI => n58, SUM(5) => N3572, SUM(4) => 
                           N3571, SUM(3) => N3570, SUM(2) => N3569, SUM(1) => 
                           N3568, SUM(0) => N3567, CO => n_1506);
   r2966 : window_rf_M4_N4_F4_NBIT32_DW01_sub_3 port map( A(31) => CWP_31_port,
                           A(30) => CWP_30_port, A(29) => CWP_29_port, A(28) =>
                           CWP_28_port, A(27) => CWP_27_port, A(26) => 
                           CWP_26_port, A(25) => CWP_25_port, A(24) => 
                           CWP_24_port, A(23) => CWP_23_port, A(22) => 
                           CWP_22_port, A(21) => CWP_21_port, A(20) => 
                           CWP_20_port, A(19) => CWP_19_port, A(18) => 
                           CWP_18_port, A(17) => CWP_17_port, A(16) => 
                           CWP_16_port, A(15) => CWP_15_port, A(14) => 
                           CWP_14_port, A(13) => CWP_13_port, A(12) => 
                           CWP_12_port, A(11) => CWP_11_port, A(10) => 
                           CWP_10_port, A(9) => CWP_9_port, A(8) => CWP_8_port,
                           A(7) => CWP_7_port, A(6) => CWP_6_port, A(5) => 
                           CWP_5_port, A(4) => CWP_4_port, A(3) => CWP_3_port, 
                           A(2) => CWP_2_port, A(1) => CWP_1_port, A(0) => 
                           CWP_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic1_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, CI => n61, DIFF(31) => N13862, 
                           DIFF(30) => N13861, DIFF(29) => N13860, DIFF(28) => 
                           N13859, DIFF(27) => N13858, DIFF(26) => N13857, 
                           DIFF(25) => N13856, DIFF(24) => N13855, DIFF(23) => 
                           N13854, DIFF(22) => N13853, DIFF(21) => N13852, 
                           DIFF(20) => N13851, DIFF(19) => N13850, DIFF(18) => 
                           N13849, DIFF(17) => N13848, DIFF(16) => N13847, 
                           DIFF(15) => N13846, DIFF(14) => N13845, DIFF(13) => 
                           N13844, DIFF(12) => N13843, DIFF(11) => N13842, 
                           DIFF(10) => N13841, DIFF(9) => N13840, DIFF(8) => 
                           N13839, DIFF(7) => N13838, DIFF(6) => N13837, 
                           DIFF(5) => N13836, DIFF(4) => N13835, DIFF(3) => 
                           N13834, DIFF(2) => N13833, DIFF(1) => N13832, 
                           DIFF(0) => N13831, CO => n_1507);
   sub_201 : window_rf_M4_N4_F4_NBIT32_DW01_sub_4 port map( A(31) => 
                           SWP_31_port, A(30) => SWP_30_port, A(29) => 
                           SWP_29_port, A(28) => SWP_28_port, A(27) => 
                           SWP_27_port, A(26) => SWP_26_port, A(25) => 
                           SWP_25_port, A(24) => SWP_24_port, A(23) => 
                           SWP_23_port, A(22) => SWP_22_port, A(21) => 
                           SWP_21_port, A(20) => SWP_20_port, A(19) => 
                           SWP_19_port, A(18) => SWP_18_port, A(17) => 
                           SWP_17_port, A(16) => SWP_16_port, A(15) => 
                           SWP_15_port, A(14) => SWP_14_port, A(13) => 
                           SWP_13_port, A(12) => SWP_12_port, A(11) => 
                           SWP_11_port, A(10) => SWP_10_port, A(9) => 
                           SWP_9_port, A(8) => SWP_8_port, A(7) => SWP_7_port, 
                           A(6) => SWP_6_port, A(5) => n846, A(4) => n841, A(3)
                           => n302, A(2) => n301, A(1) => n814, A(0) => n754, 
                           B(31) => X_Logic0_port, B(30) => X_Logic0_port, 
                           B(29) => X_Logic0_port, B(28) => X_Logic0_port, 
                           B(27) => X_Logic0_port, B(26) => X_Logic0_port, 
                           B(25) => X_Logic0_port, B(24) => X_Logic0_port, 
                           B(23) => X_Logic0_port, B(22) => X_Logic0_port, 
                           B(21) => X_Logic0_port, B(20) => X_Logic0_port, 
                           B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
                           B(17) => X_Logic0_port, B(16) => X_Logic0_port, 
                           B(15) => X_Logic0_port, B(14) => X_Logic0_port, 
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic1_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, CI => n62, 
                           DIFF(31) => N50368, DIFF(30) => N50367, DIFF(29) => 
                           N50366, DIFF(28) => N50365, DIFF(27) => N50364, 
                           DIFF(26) => N50363, DIFF(25) => N50362, DIFF(24) => 
                           N50361, DIFF(23) => N50360, DIFF(22) => N50359, 
                           DIFF(21) => N50358, DIFF(20) => N50357, DIFF(19) => 
                           N50356, DIFF(18) => N50355, DIFF(17) => N50354, 
                           DIFF(16) => N50353, DIFF(15) => N50352, DIFF(14) => 
                           N50351, DIFF(13) => N50350, DIFF(12) => N50349, 
                           DIFF(11) => N50348, DIFF(10) => N50347, DIFF(9) => 
                           N50346, DIFF(8) => N50345, DIFF(7) => N50344, 
                           DIFF(6) => N50343, DIFF(5) => N50342, DIFF(4) => 
                           N50341, DIFF(3) => N50340, DIFF(2) => n_1508, 
                           DIFF(1) => N50338, DIFF(0) => N50337, CO => n_1509);
   r2840 : window_rf_M4_N4_F4_NBIT32_DW01_add_4 port map( A(31) => CWP_31_port,
                           A(30) => CWP_30_port, A(29) => CWP_29_port, A(28) =>
                           CWP_28_port, A(27) => CWP_27_port, A(26) => 
                           CWP_26_port, A(25) => CWP_25_port, A(24) => 
                           CWP_24_port, A(23) => CWP_23_port, A(22) => 
                           CWP_22_port, A(21) => CWP_21_port, A(20) => 
                           CWP_20_port, A(19) => CWP_19_port, A(18) => 
                           CWP_18_port, A(17) => CWP_17_port, A(16) => 
                           CWP_16_port, A(15) => CWP_15_port, A(14) => 
                           CWP_14_port, A(13) => CWP_13_port, A(12) => 
                           CWP_12_port, A(11) => CWP_11_port, A(10) => 
                           CWP_10_port, A(9) => CWP_9_port, A(8) => CWP_8_port,
                           A(7) => CWP_7_port, A(6) => CWP_6_port, A(5) => 
                           CWP_5_port, A(4) => CWP_4_port, A(3) => CWP_3_port, 
                           A(2) => CWP_2_port, A(1) => CWP_1_port, A(0) => 
                           CWP_0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic1_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, CI => n65, SUM(31) => N12300, SUM(30)
                           => N12299, SUM(29) => N12298, SUM(28) => N12297, 
                           SUM(27) => N12296, SUM(26) => N12295, SUM(25) => 
                           N12294, SUM(24) => N12293, SUM(23) => N12292, 
                           SUM(22) => N12291, SUM(21) => N12290, SUM(20) => 
                           N12289, SUM(19) => N12288, SUM(18) => N12287, 
                           SUM(17) => N12286, SUM(16) => N12285, SUM(15) => 
                           N12284, SUM(14) => N12283, SUM(13) => N12282, 
                           SUM(12) => N12281, SUM(11) => N12280, SUM(10) => 
                           N12279, SUM(9) => N12278, SUM(8) => N12277, SUM(7) 
                           => N12276, SUM(6) => N12275, SUM(5) => N12274, 
                           SUM(4) => N12273, SUM(3) => N12272, SUM(2) => N12271
                           , SUM(1) => N12270, SUM(0) => N12269, CO => n_1510);
   MEM_OUT_tri_30_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_30_port);
   MEM_OUT_tri_31_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_31_port);
   MEM_OUT_tri_0_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_0_port);
   MEM_OUT_tri_1_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_1_port);
   MEM_OUT_tri_2_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_2_port);
   MEM_OUT_tri_3_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_3_port);
   MEM_OUT_tri_4_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_4_port);
   MEM_OUT_tri_5_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_5_port);
   MEM_OUT_tri_6_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_6_port);
   MEM_OUT_tri_7_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_7_port);
   MEM_OUT_tri_8_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_8_port);
   MEM_OUT_tri_9_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_9_port);
   MEM_OUT_tri_10_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_10_port);
   MEM_OUT_tri_11_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_11_port);
   MEM_OUT_tri_12_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_12_port);
   MEM_OUT_tri_13_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_13_port);
   MEM_OUT_tri_14_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_14_port);
   MEM_OUT_tri_15_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_15_port);
   MEM_OUT_tri_16_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_16_port);
   MEM_OUT_tri_17_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_17_port);
   MEM_OUT_tri_18_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_18_port);
   MEM_OUT_tri_19_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_19_port);
   MEM_OUT_tri_20_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_20_port);
   MEM_OUT_tri_21_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_21_port);
   MEM_OUT_tri_22_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_22_port);
   MEM_OUT_tri_23_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_23_port);
   MEM_OUT_tri_24_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_24_port);
   MEM_OUT_tri_25_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_25_port);
   MEM_OUT_tri_26_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_26_port);
   MEM_OUT_tri_27_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_27_port);
   MEM_OUT_tri_28_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_28_port);
   MEM_OUT_tri_29_inst : TBUF_X1 port map( A => n89, EN => n90, Z => 
                           MEM_OUT_29_port);
   SWP_reg_3_inst : DFF_X1 port map( D => n13155, CK => n977, Q => SWP_3_port, 
                           QN => n11866);
   U4 : OR2_X1 port map( A1 => n4846, A2 => n116, ZN => n2);
   U5 : OR2_X1 port map( A1 => n4809, A2 => n209, ZN => n3);
   U6 : OR3_X1 port map( A1 => n4784, A2 => n4812, A3 => n209, ZN => n4);
   U7 : OR2_X1 port map( A1 => n5183, A2 => n5184, ZN => n5);
   U8 : OR2_X1 port map( A1 => n5755, A2 => n5758, ZN => n6);
   U9 : OR2_X1 port map( A1 => n5367, A2 => n5758, ZN => n7);
   U10 : OR2_X1 port map( A1 => n6216, A2 => n6215, ZN => n8);
   U11 : OR2_X1 port map( A1 => n5755, A2 => n6215, ZN => n9);
   U12 : OR2_X1 port map( A1 => n6815, A2 => n6812, ZN => n10);
   U13 : OR3_X1 port map( A1 => n5925, A2 => n6812, A3 => n6816, ZN => n11);
   U14 : OR2_X1 port map( A1 => n7698, A2 => n7695, ZN => n12);
   U15 : OR3_X1 port map( A1 => n6823, A2 => n7695, A3 => n7699, ZN => n13);
   U16 : OR2_X1 port map( A1 => n8144, A2 => n8145, ZN => n14);
   U17 : OR3_X1 port map( A1 => n7266, A2 => n8145, A3 => n8147, ZN => n15);
   U18 : OR2_X1 port map( A1 => n8586, A2 => n8583, ZN => n16);
   U19 : OR3_X1 port map( A1 => n7707, A2 => n8583, A3 => n8587, ZN => n17);
   U21 : OR2_X1 port map( A1 => n9033, A2 => n9034, ZN => n18);
   U22 : OR3_X1 port map( A1 => n8155, A2 => n9034, A3 => n9036, ZN => n19);
   U24 : OR2_X1 port map( A1 => n9475, A2 => n9472, ZN => n20);
   U25 : OR3_X1 port map( A1 => n8596, A2 => n9472, A3 => n9476, ZN => n21);
   U27 : OR3_X1 port map( A1 => n9045, A2 => n9920, A3 => n9921, ZN => n22);
   U28 : OR2_X1 port map( A1 => n11849, A2 => n11846, ZN => n23);
   U30 : OR3_X1 port map( A1 => n9484, A2 => n11846, A3 => n11850, ZN => n24);
   U31 : OR3_X1 port map( A1 => n13489, A2 => n13631, A3 => n13632, ZN => n25);
   U34 : OR2_X1 port map( A1 => n16213, A2 => n16232, ZN => n26);
   U35 : OR2_X1 port map( A1 => n6959, A2 => n6960, ZN => n27);
   U37 : OR2_X1 port map( A1 => n7256, A2 => n7257, ZN => n28);
   U38 : OR2_X1 port map( A1 => n7402, A2 => n7403, ZN => n29);
   U39 : OR2_X1 port map( A1 => n7549, A2 => n7550, ZN => n30);
   U40 : OR2_X1 port map( A1 => n7693, A2 => n7694, ZN => n31);
   U41 : OR2_X1 port map( A1 => n7844, A2 => n7845, ZN => n32);
   U42 : OR2_X1 port map( A1 => n8140, A2 => n8141, ZN => n33);
   U43 : OR2_X1 port map( A1 => n8291, A2 => n8292, ZN => n34);
   U44 : OR2_X1 port map( A1 => n8439, A2 => n8440, ZN => n35);
   U45 : OR2_X1 port map( A1 => n8581, A2 => n8582, ZN => n36);
   U46 : OR2_X1 port map( A1 => n8732, A2 => n8733, ZN => n37);
   U47 : OR2_X1 port map( A1 => n8881, A2 => n8882, ZN => n38);
   U48 : OR2_X1 port map( A1 => n9029, A2 => n9030, ZN => n39);
   U49 : OR2_X1 port map( A1 => n9181, A2 => n9182, ZN => n40);
   U50 : OR2_X1 port map( A1 => n9328, A2 => n9329, ZN => n41);
   U51 : OR2_X1 port map( A1 => n9470, A2 => n9471, ZN => n42);
   U52 : OR2_X1 port map( A1 => n9620, A2 => n9621, ZN => n43);
   U53 : OR2_X1 port map( A1 => n9767, A2 => n9768, ZN => n44);
   U54 : OR2_X1 port map( A1 => n9914, A2 => n9915, ZN => n45);
   U55 : OR2_X1 port map( A1 => n10064, A2 => n10065, ZN => n46);
   U56 : OR2_X1 port map( A1 => n10216, A2 => n10217, ZN => n47);
   U57 : OR2_X1 port map( A1 => n11844, A2 => n11845, ZN => n48);
   U58 : OR2_X1 port map( A1 => n13328, A2 => n13329, ZN => n50);
   U59 : OR2_X1 port map( A1 => n13477, A2 => n13478, ZN => n51);
   U60 : OR2_X1 port map( A1 => n13626, A2 => n13627, ZN => n53);
   U61 : OR2_X1 port map( A1 => n4752, A2 => n4785, ZN => n54);
   U62 : AND3_X1 port map( A1 => n247, A2 => n6809, A3 => n300, ZN => n56);
   U63 : AND3_X1 port map( A1 => n293, A2 => n6958, A3 => n300, ZN => n57);
   U64 : AND3_X1 port map( A1 => n216, A2 => n6077, A3 => n300, ZN => n59);
   U65 : AND3_X1 port map( A1 => n295, A2 => n7255, A3 => n300, ZN => n60);
   U66 : AND3_X1 port map( A1 => n297, A2 => n7401, A3 => n300, ZN => n63);
   U67 : AND3_X1 port map( A1 => n299, A2 => n7548, A3 => n300, ZN => n64);
   U68 : AND3_X1 port map( A1 => n263, A2 => n7692, A3 => n300, ZN => n66);
   U69 : AND3_X1 port map( A1 => n285, A2 => n7843, A3 => n300, ZN => n67);
   U70 : AND3_X1 port map( A1 => n218, A2 => n6972, A3 => n300, ZN => n68);
   U71 : AND3_X1 port map( A1 => n265, A2 => n8139, A3 => n300, ZN => n69);
   U72 : AND3_X1 port map( A1 => n287, A2 => n8290, A3 => n300, ZN => n70);
   U73 : AND3_X1 port map( A1 => n289, A2 => n8438, A3 => n300, ZN => n71);
   U74 : AND3_X1 port map( A1 => n267, A2 => n8580, A3 => n300, ZN => n72);
   U75 : AND3_X1 port map( A1 => n291, A2 => n8731, A3 => n300, ZN => n73);
   U76 : AND3_X1 port map( A1 => n277, A2 => n8880, A3 => n300, ZN => n74);
   U77 : AND3_X1 port map( A1 => n253, A2 => n9028, A3 => n300, ZN => n75);
   U78 : AND3_X1 port map( A1 => n279, A2 => n9180, A3 => n300, ZN => n76);
   U79 : AND3_X1 port map( A1 => n281, A2 => n9327, A3 => n300, ZN => n77);
   U80 : AND3_X1 port map( A1 => n255, A2 => n9469, A3 => n300, ZN => n78);
   U81 : AND3_X1 port map( A1 => n283, A2 => n9619, A3 => n300, ZN => n79);
   U82 : AND3_X1 port map( A1 => n269, A2 => n9766, A3 => n300, ZN => n80);
   U83 : AND3_X1 port map( A1 => n257, A2 => n9913, A3 => n300, ZN => n81);
   U84 : AND3_X1 port map( A1 => n271, A2 => n10063, A3 => n300, ZN => n82);
   U85 : AND3_X1 port map( A1 => n273, A2 => n10215, A3 => n300, ZN => n83);
   U86 : AND3_X1 port map( A1 => n259, A2 => n11843, A3 => n300, ZN => n84);
   U87 : AND3_X1 port map( A1 => n275, A2 => n13327, A3 => n300, ZN => n85);
   U88 : AND3_X1 port map( A1 => n261, A2 => n13476, A3 => n300, ZN => n86);
   U89 : AND3_X1 port map( A1 => n245, A2 => n13625, A3 => n300, ZN => n87);
   U90 : AND3_X1 port map( A1 => n249, A2 => n9927, A3 => n300, ZN => n88);
   U91 : AND3_X1 port map( A1 => n251, A2 => n10078, A3 => n300, ZN => n91);
   U92 : OR2_X1 port map( A1 => n4752, A2 => n4784, ZN => n92);
   U93 : OR2_X1 port map( A1 => n5515, A2 => n5758, ZN => n93);
   U94 : OR2_X1 port map( A1 => n5756, A2 => n5758, ZN => n94);
   U95 : OR2_X1 port map( A1 => n6066, A2 => n6215, ZN => n95);
   U96 : OR2_X1 port map( A1 => n6217, A2 => n6215, ZN => n96);
   U97 : OR2_X1 port map( A1 => n6671, A2 => n6812, ZN => n97);
   U98 : OR2_X1 port map( A1 => n6521, A2 => n6812, ZN => n98);
   U99 : OR2_X1 port map( A1 => n7553, A2 => n7695, ZN => n99);
   U100 : OR2_X1 port map( A1 => n7406, A2 => n7695, ZN => n100);
   U101 : OR2_X1 port map( A1 => n8443, A2 => n8583, ZN => n101);
   U102 : OR2_X1 port map( A1 => n8295, A2 => n8583, ZN => n102);
   U103 : OR2_X1 port map( A1 => n9332, A2 => n9472, ZN => n103);
   U104 : OR2_X1 port map( A1 => n9185, A2 => n9472, ZN => n104);
   U105 : OR2_X1 port map( A1 => n10219, A2 => n11846, ZN => n105);
   U106 : OR2_X1 port map( A1 => n10067, A2 => n11846, ZN => n106);
   U107 : OR2_X1 port map( A1 => n13781, A2 => n13782, ZN => n107);
   U108 : OR2_X1 port map( A1 => n13781, A2 => n16232, ZN => n108);
   U109 : OR2_X1 port map( A1 => n6214, A2 => n6215, ZN => n109);
   U110 : OR3_X1 port map( A1 => n6812, A2 => n6369, A3 => n6813, ZN => n110);
   U111 : OR3_X1 port map( A1 => n7695, A2 => n7261, A3 => n7696, ZN => n111);
   U112 : OR3_X1 port map( A1 => n8583, A2 => n8153, A3 => n8584, ZN => n112);
   U113 : OR3_X1 port map( A1 => n9472, A2 => n9042, A3 => n9473, ZN => n113);
   U114 : OR3_X1 port map( A1 => n11846, A2 => n9918, A3 => n11847, ZN => n114)
                           ;
   U115 : OR2_X1 port map( A1 => n2, A2 => n13796, ZN => n115);
   U116 : NOR3_X2 port map( A1 => n840, A2 => n11867, A3 => n813, ZN => n5775);
   U117 : NOR3_X2 port map( A1 => SWP_4_port, A2 => n11864, A3 => SWP_3_port, 
                           ZN => n5216);
   U118 : NOR3_X2 port map( A1 => SWP_3_port, A2 => n11865, A3 => SWP_5_port, 
                           ZN => n7708);
   U119 : NOR3_X2 port map( A1 => SWP_4_port, A2 => n11866, A3 => SWP_5_port, 
                           ZN => n8895);
   U120 : NOR3_X2 port map( A1 => SWP_3_port, A2 => SWP_4_port, A3 => 
                           SWP_5_port, ZN => n10080);
   U121 : NOR3_X2 port map( A1 => CWP_1_port, A2 => n11863, A3 => CWP_2_port, 
                           ZN => n16286);
   U122 : NOR3_X2 port map( A1 => n11865, A2 => n11866, A3 => SWP_5_port, ZN =>
                           n6531);
   U123 : INV_X1 port map( A => n13862_port, ZN => n118);
   U124 : INV_X2 port map( A => n118, ZN => n119);
   U125 : INV_X2 port map( A => n5356, ZN => n5220);
   U126 : INV_X2 port map( A => n5512, ZN => n5376);
   U127 : AND2_X2 port map( A1 => n7111, A2 => n7112, ZN => n6977);
   U128 : AND2_X2 port map( A1 => n7996, A2 => n7997, ZN => n7862);
   U129 : AND2_X2 port map( A1 => n8884, A2 => n8885, ZN => n8749);
   U130 : AND2_X2 port map( A1 => n9770, A2 => n9771, ZN => n9635);
   U131 : AND2_X2 port map( A1 => n13480, A2 => n13481, ZN => n13345);
   U132 : AND2_X2 port map( A1 => n5193, A2 => n5358, ZN => n5228);
   U133 : AND2_X2 port map( A1 => n5360, A2 => n5514, ZN => n5382);
   U134 : AND2_X2 port map( A1 => n5194, A2 => n5514, ZN => n5384);
   U135 : AND2_X2 port map( A1 => n5769, A2 => n5915, ZN => n5785);
   U136 : AND2_X2 port map( A1 => n5517, A2 => n5915, ZN => n5787);
   U137 : AND2_X2 port map( A1 => n5917, A2 => n6067, ZN => n5936);
   U138 : AND2_X2 port map( A1 => n5769, A2 => n6067, ZN => n5938);
   U139 : AND2_X2 port map( A1 => n6224, A2 => n6367, ZN => n6238);
   U140 : AND2_X2 port map( A1 => n6069, A2 => n6367, ZN => n6240);
   U141 : AND2_X2 port map( A1 => n6369, A2 => n6520, ZN => n6391);
   U142 : AND2_X2 port map( A1 => n6224, A2 => n6520, ZN => n6393);
   U143 : AND2_X2 port map( A1 => n6522, A2 => n6670, ZN => n6541);
   U144 : AND2_X2 port map( A1 => n6369, A2 => n6670, ZN => n6543);
   U145 : AND2_X2 port map( A1 => n6963, A2 => n6962, ZN => n6831);
   U146 : AND2_X2 port map( A1 => n6672, A2 => n6962, ZN => n6833);
   U147 : AND2_X2 port map( A1 => n6964, A2 => n7112, ZN => n6982);
   U148 : AND2_X2 port map( A1 => n6963, A2 => n7112, ZN => n6984);
   U149 : AND2_X2 port map( A1 => n7113, A2 => n7259, ZN => n7128);
   U150 : AND2_X2 port map( A1 => n6964, A2 => n7259, ZN => n7130);
   U151 : AND2_X2 port map( A1 => n7261, A2 => n7405, ZN => n7274);
   U152 : AND2_X2 port map( A1 => n7113, A2 => n7405, ZN => n7276);
   U153 : AND2_X2 port map( A1 => n7407, A2 => n7552, ZN => n7421);
   U154 : AND2_X2 port map( A1 => n7261, A2 => n7552, ZN => n7423);
   U155 : AND2_X2 port map( A1 => n7849, A2 => n7848, ZN => n7716);
   U156 : AND2_X2 port map( A1 => n7554, A2 => n7848, ZN => n7718);
   U157 : AND2_X2 port map( A1 => n7850, A2 => n7997, ZN => n7867);
   U158 : AND2_X2 port map( A1 => n7849, A2 => n7997, ZN => n7869);
   U159 : AND2_X2 port map( A1 => n7998, A2 => n8143, ZN => n8013);
   U160 : AND2_X2 port map( A1 => n8153, A2 => n8294, ZN => n8163);
   U161 : AND2_X2 port map( A1 => n7998, A2 => n8294, ZN => n8165);
   U162 : AND2_X2 port map( A1 => n8296, A2 => n8442, ZN => n8311);
   U163 : AND2_X2 port map( A1 => n8153, A2 => n8442, ZN => n8313);
   U164 : AND2_X2 port map( A1 => n8593, A2 => n8736, ZN => n8604);
   U165 : AND2_X2 port map( A1 => n8444, A2 => n8736, ZN => n8606);
   U166 : AND2_X2 port map( A1 => n8737, A2 => n8885, ZN => n8753);
   U167 : AND2_X2 port map( A1 => n8593, A2 => n8885, ZN => n8755);
   U168 : AND2_X2 port map( A1 => n8886, A2 => n9032, ZN => n8902);
   U169 : AND2_X2 port map( A1 => n9042, A2 => n9184, ZN => n9053);
   U170 : AND2_X2 port map( A1 => n8886, A2 => n9184, ZN => n9055);
   U171 : AND2_X2 port map( A1 => n9186, A2 => n9331, ZN => n9200);
   U172 : AND2_X2 port map( A1 => n9042, A2 => n9331, ZN => n9202);
   U173 : AND2_X2 port map( A1 => n9482, A2 => n9624, ZN => n9492);
   U174 : AND2_X2 port map( A1 => n9333, A2 => n9624, ZN => n9494);
   U175 : AND2_X2 port map( A1 => n9625, A2 => n9771, ZN => n9639);
   U176 : AND2_X2 port map( A1 => n9482, A2 => n9771, ZN => n9641);
   U177 : AND2_X2 port map( A1 => n9772, A2 => n9917, ZN => n9787);
   U178 : AND2_X2 port map( A1 => n9918, A2 => n10066, ZN => n9936);
   U179 : AND2_X2 port map( A1 => n9772, A2 => n10066, ZN => n9938);
   U180 : AND2_X2 port map( A1 => n10068, A2 => n10218, ZN => n10088);
   U181 : AND2_X2 port map( A1 => n9918, A2 => n10218, ZN => n10090);
   U182 : AND2_X2 port map( A1 => n13333, A2 => n13332, ZN => n13200);
   U183 : AND2_X2 port map( A1 => n10220, A2 => n13332, ZN => n13202);
   U184 : AND2_X2 port map( A1 => n10220, A2 => n13481, ZN => n13349);
   U185 : AND2_X2 port map( A1 => n13482, A2 => n13481, ZN => n13351);
   U186 : AND2_X2 port map( A1 => n13633, A2 => n13629, ZN => n13500);
   U187 : AND2_X2 port map( A1 => n13633, A2 => n13780, ZN => n13653);
   U188 : AND2_X2 port map( A1 => n13633, A2 => n16212, ZN => n13881);
   U189 : AND2_X2 port map( A1 => n5197, A2 => n5187, ZN => n4874);
   U190 : AND2_X2 port map( A1 => n5194, A2 => n5358, ZN => n5226);
   U191 : AND3_X2 port map( A1 => n11848, A2 => n13331, A3 => n13332, ZN => 
                           n13196);
   U192 : AND2_X2 port map( A1 => n5193, A2 => n5187, ZN => n4870);
   U193 : AND3_X2 port map( A1 => n8585, A2 => n8735, A3 => n8736, ZN => n8600)
                           ;
   U194 : AND3_X2 port map( A1 => n9474, A2 => n9623, A3 => n9624, ZN => n9488)
                           ;
   U195 : AND3_X2 port map( A1 => n6814, A2 => n6961, A3 => n6962, ZN => n6827)
                           ;
   U196 : AND3_X2 port map( A1 => n7697, A2 => n7847, A3 => n7848, ZN => n7712)
                           ;
   U197 : AND3_X2 port map( A1 => n5915, A2 => n5756, A3 => n5916, ZN => n5779)
                           ;
   U198 : AND3_X2 port map( A1 => n5916, A2 => n6066, A3 => n6067, ZN => n5930)
                           ;
   U199 : AND4_X2 port map( A1 => n16212, A2 => n13628, A3 => n16213, A4 => 
                           n13781, ZN => n13792);
   U200 : AND3_X2 port map( A1 => n5762, A2 => n5763, A3 => n300, ZN => n5530);
   U201 : AND4_X2 port map( A1 => n10066, A2 => n9916, A3 => n9623, A4 => 
                           n10067, ZN => n9932);
   U202 : AND4_X2 port map( A1 => n10218, A2 => n9916, A3 => n10067, A4 => 
                           n10219, ZN => n10084);
   U203 : AND4_X2 port map( A1 => n9184, A2 => n9031, A3 => n8735, A4 => n9185,
                           ZN => n9049);
   U204 : AND4_X2 port map( A1 => n9331, A2 => n9031, A3 => n9185, A4 => n9332,
                           ZN => n9196);
   U205 : AND4_X2 port map( A1 => n8294, A2 => n8142, A3 => n7847, A4 => n8295,
                           ZN => n8159);
   U206 : AND4_X2 port map( A1 => n8442, A2 => n8142, A3 => n8295, A4 => n8443,
                           ZN => n8307);
   U207 : AND4_X2 port map( A1 => n7405, A2 => n7260, A3 => n6961, A4 => n7406,
                           ZN => n7270);
   U208 : AND4_X2 port map( A1 => n7552, A2 => n7260, A3 => n7406, A4 => n7553,
                           ZN => n7417);
   U209 : AND4_X2 port map( A1 => n6670, A2 => n6368, A3 => n6521, A4 => n6671,
                           ZN => n6535);
   U210 : AND4_X2 port map( A1 => n7259, A2 => n7260, A3 => n6815, A4 => n6961,
                           ZN => n7124);
   U211 : AND4_X2 port map( A1 => n6367, A2 => n6368, A3 => n6217, A4 => n6066,
                           ZN => n6232);
   U212 : AND4_X2 port map( A1 => n6520, A2 => n6368, A3 => n6066, A4 => n6521,
                           ZN => n6385);
   U213 : AND2_X2 port map( A1 => n16210, A2 => n16211, ZN => n13793);
   U214 : INV_X2 port map( A => n5185, ZN => n4862);
   U215 : AND2_X2 port map( A1 => n6810, A2 => n6811, ZN => n6682);
   U216 : AND2_X2 port map( A1 => n13778, A2 => n13779, ZN => n13648);
   U217 : INV_X2 port map( A => n88, ZN => n120);
   U218 : INV_X2 port map( A => n91, ZN => n121);
   U219 : INV_X2 port map( A => n86, ZN => n122);
   U220 : INV_X2 port map( A => n87, ZN => n123);
   U221 : INV_X2 port map( A => n84, ZN => n124);
   U222 : INV_X2 port map( A => n85, ZN => n125);
   U223 : INV_X2 port map( A => n82, ZN => n126);
   U224 : INV_X2 port map( A => n83, ZN => n127);
   U225 : INV_X2 port map( A => n80, ZN => n128);
   U226 : INV_X2 port map( A => n81, ZN => n129);
   U227 : INV_X2 port map( A => n78, ZN => n130);
   U228 : INV_X2 port map( A => n79, ZN => n131);
   U229 : INV_X2 port map( A => n76, ZN => n132);
   U230 : INV_X2 port map( A => n77, ZN => n133);
   U231 : INV_X2 port map( A => n74, ZN => n134);
   U232 : INV_X2 port map( A => n75, ZN => n135);
   U233 : INV_X2 port map( A => n72, ZN => n136);
   U234 : INV_X2 port map( A => n73, ZN => n137);
   U235 : INV_X2 port map( A => n70, ZN => n138);
   U236 : INV_X2 port map( A => n71, ZN => n139);
   U237 : INV_X2 port map( A => n68, ZN => n140);
   U238 : INV_X2 port map( A => n69, ZN => n141);
   U239 : INV_X2 port map( A => n66, ZN => n142);
   U240 : INV_X2 port map( A => n67, ZN => n143);
   U241 : INV_X2 port map( A => n63, ZN => n144);
   U242 : INV_X2 port map( A => n64, ZN => n145);
   U243 : INV_X2 port map( A => n59, ZN => n146);
   U244 : INV_X2 port map( A => n60, ZN => n147);
   U245 : INV_X2 port map( A => n56, ZN => n148);
   U246 : INV_X2 port map( A => n57, ZN => n149);
   U247 : NAND3_X2 port map( A1 => n226, A2 => n5370, A3 => n300, ZN => n6389);
   U248 : NAND3_X2 port map( A1 => n228, A2 => n5524, A3 => n300, ZN => n6539);
   U249 : NAND3_X2 port map( A1 => n6085, A2 => n6211, A3 => n300, ZN => n6086)
                           ;
   U250 : NAND3_X2 port map( A1 => n224, A2 => n5213, A3 => n300, ZN => n6236);
   U251 : NAND3_X2 port map( A1 => n235, A2 => n5912, A3 => n300, ZN => n5783);
   U252 : NAND3_X2 port map( A1 => n222, A2 => n6063, A3 => n300, ZN => n5934);
   U253 : NAND3_X2 port map( A1 => n231, A2 => n5353, A3 => n300, ZN => n5224);
   U254 : NAND3_X2 port map( A1 => n233, A2 => n5509, A3 => n300, ZN => n5380);
   U255 : AND2_X2 port map( A1 => n13482, A2 => n13780, ZN => n13652);
   U256 : AND2_X2 port map( A1 => n13482, A2 => n16212, ZN => n13880);
   U257 : AND2_X2 port map( A1 => n13333, A2 => n13481, ZN => n13350);
   U258 : AND2_X2 port map( A1 => n13482, A2 => n13629, ZN => n13499);
   U259 : AND2_X2 port map( A1 => n10068, A2 => n13332, ZN => n13201);
   U260 : AND2_X2 port map( A1 => n13334, A2 => n13481, ZN => n13348);
   U261 : AND2_X2 port map( A1 => n9772, A2 => n10218, ZN => n10089);
   U262 : AND2_X2 port map( A1 => n13334, A2 => n13332, ZN => n13199);
   U263 : AND2_X2 port map( A1 => n9919, A2 => n10066, ZN => n9937);
   U264 : AND2_X2 port map( A1 => n10220, A2 => n10218, ZN => n10087);
   U265 : AND2_X2 port map( A1 => n9918, A2 => n9917, ZN => n9786);
   U266 : AND2_X2 port map( A1 => n10068, A2 => n10066, ZN => n9935);
   U267 : AND2_X2 port map( A1 => n9772, A2 => n9771, ZN => n9638);
   U268 : AND2_X2 port map( A1 => n9333, A2 => n9771, ZN => n9640);
   U269 : AND2_X2 port map( A1 => n9625, A2 => n9624, ZN => n9491);
   U270 : AND2_X2 port map( A1 => n9186, A2 => n9624, ZN => n9493);
   U271 : AND2_X2 port map( A1 => n9333, A2 => n9331, ZN => n9199);
   U272 : AND2_X2 port map( A1 => n8886, A2 => n9331, ZN => n9201);
   U273 : AND2_X2 port map( A1 => n9186, A2 => n9184, ZN => n9052);
   U274 : AND2_X2 port map( A1 => n9035, A2 => n9184, ZN => n9054);
   U275 : AND2_X2 port map( A1 => n8886, A2 => n8885, ZN => n8752);
   U276 : AND2_X2 port map( A1 => n8444, A2 => n8885, ZN => n8754);
   U277 : AND2_X2 port map( A1 => n8737, A2 => n8736, ZN => n8603);
   U278 : AND2_X2 port map( A1 => n8296, A2 => n8736, ZN => n8605);
   U279 : AND2_X2 port map( A1 => n8444, A2 => n8442, ZN => n8310);
   U280 : AND2_X2 port map( A1 => n7998, A2 => n8442, ZN => n8312);
   U281 : AND2_X2 port map( A1 => n8296, A2 => n8294, ZN => n8162);
   U282 : AND2_X2 port map( A1 => n8146, A2 => n8294, ZN => n8164);
   U283 : AND2_X2 port map( A1 => n7998, A2 => n7997, ZN => n7866);
   U284 : AND2_X2 port map( A1 => n7554, A2 => n7997, ZN => n7868);
   U285 : AND2_X2 port map( A1 => n7850, A2 => n7848, ZN => n7715);
   U286 : AND2_X2 port map( A1 => n7407, A2 => n7848, ZN => n7717);
   U287 : AND2_X2 port map( A1 => n7554, A2 => n7552, ZN => n7420);
   U288 : AND2_X2 port map( A1 => n7113, A2 => n7552, ZN => n7422);
   U289 : AND2_X2 port map( A1 => n7407, A2 => n7405, ZN => n7273);
   U290 : AND2_X2 port map( A1 => n6964, A2 => n7405, ZN => n7275);
   U291 : AND2_X2 port map( A1 => n7261, A2 => n7259, ZN => n7127);
   U292 : AND2_X2 port map( A1 => n6963, A2 => n7259, ZN => n7129);
   U293 : AND2_X2 port map( A1 => n7113, A2 => n7112, ZN => n6981);
   U294 : AND2_X2 port map( A1 => n6672, A2 => n7112, ZN => n6983);
   U295 : AND2_X2 port map( A1 => n6964, A2 => n6962, ZN => n6830);
   U296 : AND2_X2 port map( A1 => n6522, A2 => n6962, ZN => n6832);
   U297 : AND2_X2 port map( A1 => n6672, A2 => n6670, ZN => n6540);
   U298 : AND2_X2 port map( A1 => n6224, A2 => n6670, ZN => n6542);
   U299 : AND2_X2 port map( A1 => n6522, A2 => n6520, ZN => n6390);
   U300 : AND2_X2 port map( A1 => n6069, A2 => n6520, ZN => n6392);
   U301 : AND2_X2 port map( A1 => n6369, A2 => n6367, ZN => n6237);
   U302 : AND2_X2 port map( A1 => n5917, A2 => n6367, ZN => n6239);
   U303 : AND2_X2 port map( A1 => n6069, A2 => n6067, ZN => n5935);
   U304 : AND2_X2 port map( A1 => n5517, A2 => n6067, ZN => n5937);
   U305 : AND2_X2 port map( A1 => n5193, A2 => n5514, ZN => n5383);
   U306 : AND2_X2 port map( A1 => n5917, A2 => n5915, ZN => n5784);
   U307 : AND2_X2 port map( A1 => n5197, A2 => n5358, ZN => n5227);
   U308 : AND2_X2 port map( A1 => n5517, A2 => n5514, ZN => n5381);
   U309 : AND2_X2 port map( A1 => n5194, A2 => n5187, ZN => n4868);
   U310 : AND2_X2 port map( A1 => n5360, A2 => n5358, ZN => n5225);
   U311 : AND3_X2 port map( A1 => n5359, A2 => n5915, A3 => n5918, ZN => n5786)
                           ;
   U312 : AND3_X2 port map( A1 => n5189, A2 => n5187, A3 => n5198, ZN => n4872)
                           ;
   U313 : NAND3_X2 port map( A1 => n4865, A2 => n5182, A3 => n300, ZN => n4866)
                           ;
   U314 : INV_X2 port map( A => n5762, ZN => n5532);
   U315 : NAND2_X2 port map( A1 => ENABLE, A2 => n16346, ZN => n4752);
   U316 : NAND4_X2 port map( A1 => n5515, A2 => n5755, A3 => n5756, A4 => n5757
                           , ZN => n5537);
   U317 : NAND2_X2 port map( A1 => n16170, A2 => n16171, ZN => n5175);
   U318 : NAND2_X2 port map( A1 => n16094, A2 => n16095, ZN => n5165);
   U319 : NAND2_X2 port map( A1 => n16134, A2 => n16135, ZN => n5173);
   U320 : NAND2_X2 port map( A1 => n15982, A2 => n15983, ZN => n5153);
   U321 : NAND2_X2 port map( A1 => n16018, A2 => n16019, ZN => n5155);
   U322 : NAND2_X2 port map( A1 => n15790, A2 => n15791, ZN => n5125);
   U323 : NAND2_X2 port map( A1 => n15942, A2 => n15943, ZN => n5145);
   U324 : NAND2_X2 port map( A1 => n15714, A2 => n15715, ZN => n5115);
   U325 : NAND2_X2 port map( A1 => n15754, A2 => n15755, ZN => n5123);
   U326 : NAND2_X2 port map( A1 => n15526, A2 => n15527, ZN => n5093);
   U327 : NAND2_X2 port map( A1 => n15562, A2 => n15563, ZN => n5095);
   U328 : NAND2_X2 port map( A1 => n15334, A2 => n15335, ZN => n5065);
   U329 : NAND2_X2 port map( A1 => n15486, A2 => n15487, ZN => n5085);
   U330 : NAND2_X2 port map( A1 => n15258, A2 => n15259, ZN => n5055);
   U331 : NAND2_X2 port map( A1 => n15298, A2 => n15299, ZN => n5063);
   U332 : NAND2_X2 port map( A1 => n15070, A2 => n15071, ZN => n5033);
   U333 : NAND2_X2 port map( A1 => n15106, A2 => n15107, ZN => n5035);
   U334 : NAND2_X2 port map( A1 => n14878, A2 => n14879, ZN => n5005);
   U335 : NAND2_X2 port map( A1 => n15030, A2 => n15031, ZN => n5025);
   U336 : NAND2_X2 port map( A1 => n14802, A2 => n14803, ZN => n4995);
   U337 : NAND2_X2 port map( A1 => n14842, A2 => n14843, ZN => n5003);
   U338 : NAND2_X2 port map( A1 => n14614, A2 => n14615, ZN => n4973);
   U339 : NAND2_X2 port map( A1 => n14650, A2 => n14651, ZN => n4975);
   U340 : NAND2_X2 port map( A1 => n14422, A2 => n14423, ZN => n4945);
   U341 : NAND2_X2 port map( A1 => n14574, A2 => n14575, ZN => n4965);
   U342 : NAND2_X2 port map( A1 => n14346, A2 => n14347, ZN => n4935);
   U343 : NAND2_X2 port map( A1 => n14386, A2 => n14387, ZN => n4943);
   U344 : NAND2_X2 port map( A1 => n14158, A2 => n14159, ZN => n4913);
   U345 : NAND2_X2 port map( A1 => n14194, A2 => n14195, ZN => n4915);
   U346 : NAND2_X2 port map( A1 => n14118, A2 => n14119, ZN => n4905);
   U347 : INV_X2 port map( A => n108, ZN => n150);
   U348 : INV_X2 port map( A => n109, ZN => n151);
   U349 : INV_X2 port map( A => n106, ZN => n152);
   U350 : INV_X2 port map( A => n107, ZN => n153);
   U351 : INV_X2 port map( A => n104, ZN => n154);
   U352 : INV_X2 port map( A => n105, ZN => n155);
   U353 : INV_X2 port map( A => n102, ZN => n156);
   U354 : INV_X2 port map( A => n103, ZN => n157);
   U355 : INV_X2 port map( A => n100, ZN => n158);
   U356 : INV_X2 port map( A => n101, ZN => n159);
   U357 : INV_X2 port map( A => n98, ZN => n160);
   U358 : INV_X2 port map( A => n99, ZN => n161);
   U359 : INV_X2 port map( A => n96, ZN => n162);
   U360 : INV_X2 port map( A => n97, ZN => n163);
   U361 : INV_X2 port map( A => n94, ZN => n164);
   U362 : INV_X2 port map( A => n95, ZN => n165);
   U363 : INV_X2 port map( A => n92, ZN => n166);
   U364 : INV_X2 port map( A => n93, ZN => n167);
   U365 : INV_X2 port map( A => n53, ZN => n168);
   U366 : INV_X2 port map( A => n54, ZN => n169);
   U367 : INV_X2 port map( A => n50, ZN => n170);
   U368 : INV_X2 port map( A => n51, ZN => n171);
   U369 : INV_X2 port map( A => n47, ZN => n172);
   U370 : INV_X2 port map( A => n48, ZN => n173);
   U371 : INV_X2 port map( A => n45, ZN => n174);
   U372 : INV_X2 port map( A => n46, ZN => n175);
   U373 : INV_X2 port map( A => n43, ZN => n176);
   U374 : INV_X2 port map( A => n44, ZN => n177);
   U375 : INV_X2 port map( A => n39, ZN => n178);
   U376 : INV_X2 port map( A => n40, ZN => n179);
   U377 : INV_X2 port map( A => n41, ZN => n180);
   U378 : INV_X2 port map( A => n42, ZN => n181);
   U379 : INV_X2 port map( A => n35, ZN => n182);
   U380 : INV_X2 port map( A => n36, ZN => n183);
   U381 : INV_X2 port map( A => n37, ZN => n184);
   U382 : INV_X2 port map( A => n38, ZN => n185);
   U383 : INV_X2 port map( A => n31, ZN => n186);
   U384 : INV_X2 port map( A => n32, ZN => n187);
   U385 : INV_X2 port map( A => n33, ZN => n188);
   U386 : INV_X2 port map( A => n34, ZN => n189);
   U387 : INV_X2 port map( A => n27, ZN => n190);
   U388 : INV_X2 port map( A => n28, ZN => n191);
   U389 : INV_X2 port map( A => n29, ZN => n192);
   U390 : INV_X2 port map( A => n30, ZN => n193);
   U391 : INV_X2 port map( A => n18, ZN => n194);
   U392 : INV_X2 port map( A => n20, ZN => n195);
   U393 : INV_X2 port map( A => n23, ZN => n196);
   U394 : INV_X2 port map( A => n26, ZN => n197);
   U395 : INV_X2 port map( A => n10, ZN => n198);
   U396 : INV_X2 port map( A => n12, ZN => n199);
   U397 : INV_X2 port map( A => n14, ZN => n200);
   U398 : INV_X2 port map( A => n16, ZN => n201);
   U399 : INV_X2 port map( A => n6, ZN => n202);
   U400 : INV_X2 port map( A => n7, ZN => n203);
   U401 : INV_X2 port map( A => n8, ZN => n204);
   U402 : INV_X2 port map( A => n9, ZN => n205);
   U403 : INV_X2 port map( A => n5, ZN => n206);
   U404 : INV_X2 port map( A => n3, ZN => n207);
   U405 : INV_X4 port map( A => n115, ZN => n208);
   U406 : INV_X1 port map( A => n4851, ZN => n209);
   U407 : INV_X2 port map( A => n209, ZN => n210);
   U408 : INV_X2 port map( A => n112, ZN => n211);
   U409 : INV_X2 port map( A => n113, ZN => n212);
   U410 : INV_X2 port map( A => n114, ZN => n213);
   U411 : INV_X2 port map( A => n4, ZN => n214);
   U412 : INV_X1 port map( A => n6980, ZN => n215);
   U413 : INV_X2 port map( A => n215, ZN => n216);
   U414 : INV_X1 port map( A => n7865, ZN => n217);
   U415 : INV_X2 port map( A => n217, ZN => n218);
   U416 : INV_X2 port map( A => n110, ZN => n219);
   U417 : INV_X2 port map( A => n111, ZN => n220);
   U418 : INV_X1 port map( A => n5933, ZN => n221);
   U419 : INV_X2 port map( A => n221, ZN => n222);
   U420 : INV_X1 port map( A => n6235, ZN => n223);
   U421 : INV_X2 port map( A => n223, ZN => n224);
   U422 : INV_X1 port map( A => n6388, ZN => n225);
   U423 : INV_X2 port map( A => n225, ZN => n226);
   U424 : INV_X1 port map( A => n6538, ZN => n227);
   U425 : INV_X2 port map( A => n227, ZN => n228);
   U426 : INV_X2 port map( A => n25, ZN => n229);
   U427 : INV_X1 port map( A => n5223, ZN => n230);
   U428 : INV_X2 port map( A => n230, ZN => n231);
   U429 : INV_X1 port map( A => n5379, ZN => n232);
   U430 : INV_X2 port map( A => n232, ZN => n233);
   U431 : INV_X1 port map( A => n5782, ZN => n234);
   U432 : INV_X2 port map( A => n234, ZN => n235);
   U433 : INV_X2 port map( A => n19, ZN => n236);
   U434 : INV_X2 port map( A => n21, ZN => n237);
   U435 : INV_X2 port map( A => n22, ZN => n238);
   U436 : INV_X2 port map( A => n24, ZN => n239);
   U437 : INV_X2 port map( A => n11, ZN => n240);
   U438 : INV_X2 port map( A => n13, ZN => n241);
   U439 : INV_X2 port map( A => n15, ZN => n242);
   U440 : INV_X2 port map( A => n17, ZN => n243);
   U441 : INV_X1 port map( A => n13497, ZN => n244);
   U442 : INV_X2 port map( A => n244, ZN => n245);
   U443 : INV_X1 port map( A => n6684, ZN => n246);
   U444 : INV_X2 port map( A => n246, ZN => n247);
   U445 : INV_X1 port map( A => n13650, ZN => n248);
   U446 : INV_X2 port map( A => n248, ZN => n249);
   U447 : INV_X1 port map( A => n13795, ZN => n250);
   U448 : INV_X2 port map( A => n250, ZN => n251);
   U449 : INV_X1 port map( A => n8901, ZN => n252);
   U450 : INV_X2 port map( A => n252, ZN => n253);
   U451 : INV_X1 port map( A => n9344, ZN => n254);
   U452 : INV_X2 port map( A => n254, ZN => n255);
   U453 : INV_X1 port map( A => n9785, ZN => n256);
   U454 : INV_X2 port map( A => n256, ZN => n257);
   U455 : INV_X1 port map( A => n10231, ZN => n258);
   U456 : INV_X2 port map( A => n258, ZN => n259);
   U457 : INV_X1 port map( A => n13347, ZN => n260);
   U458 : INV_X2 port map( A => n260, ZN => n261);
   U459 : INV_X1 port map( A => n7567, ZN => n262);
   U460 : INV_X2 port map( A => n262, ZN => n263);
   U461 : INV_X1 port map( A => n8012, ZN => n264);
   U462 : INV_X2 port map( A => n264, ZN => n265);
   U463 : INV_X1 port map( A => n8455, ZN => n266);
   U464 : INV_X2 port map( A => n266, ZN => n267);
   U465 : INV_X1 port map( A => n9637, ZN => n268);
   U466 : INV_X2 port map( A => n268, ZN => n269);
   U467 : INV_X1 port map( A => n9934, ZN => n270);
   U468 : INV_X2 port map( A => n270, ZN => n271);
   U469 : INV_X1 port map( A => n10086, ZN => n272);
   U470 : INV_X2 port map( A => n272, ZN => n273);
   U471 : INV_X1 port map( A => n13198, ZN => n274);
   U472 : INV_X2 port map( A => n274, ZN => n275);
   U473 : INV_X1 port map( A => n8751, ZN => n276);
   U474 : INV_X2 port map( A => n276, ZN => n277);
   U475 : INV_X1 port map( A => n9051, ZN => n278);
   U476 : INV_X2 port map( A => n278, ZN => n279);
   U477 : INV_X1 port map( A => n9198, ZN => n280);
   U478 : INV_X2 port map( A => n280, ZN => n281);
   U479 : INV_X1 port map( A => n9490, ZN => n282);
   U480 : INV_X2 port map( A => n282, ZN => n283);
   U481 : INV_X1 port map( A => n7714, ZN => n284);
   U482 : INV_X2 port map( A => n284, ZN => n285);
   U483 : INV_X1 port map( A => n8161, ZN => n286);
   U484 : INV_X2 port map( A => n286, ZN => n287);
   U485 : INV_X1 port map( A => n8309, ZN => n288);
   U486 : INV_X2 port map( A => n288, ZN => n289);
   U487 : INV_X1 port map( A => n8602, ZN => n290);
   U488 : INV_X2 port map( A => n290, ZN => n291);
   U489 : INV_X1 port map( A => n6829, ZN => n292);
   U490 : INV_X2 port map( A => n292, ZN => n293);
   U491 : INV_X1 port map( A => n7126, ZN => n294);
   U492 : INV_X2 port map( A => n294, ZN => n295);
   U493 : INV_X1 port map( A => n7272, ZN => n296);
   U494 : INV_X2 port map( A => n296, ZN => n297);
   U495 : INV_X1 port map( A => n7419, ZN => n298);
   U496 : INV_X2 port map( A => n298, ZN => n299);
   U497 : OAI221_X4 port map( B1 => n4786, B2 => n5202, C1 => n5203, C2 => 
                           n5204, A => n5205, ZN => n4865);
   U498 : OAI22_X4 port map( A1 => n4786, A2 => n6220, B1 => n6221, B2 => n5204
                           , ZN => n6085);
   U499 : OAI21_X4 port map( B1 => n4788, B2 => n4812, A => ENABLE, ZN => n5204
                           );
   U500 : INV_X2 port map( A => n2, ZN => n300);
   U501 : INV_X4 port map( A => n5206, ZN => n4787);
   U502 : NOR2_X4 port map( A1 => n4840, A2 => n4785, ZN => n5206);
   U503 : AND2_X4 port map( A1 => n16243, A2 => n16244, ZN => n13825);
   U504 : INV_X4 port map( A => n13890, ZN => n13807);
   U505 : AND2_X4 port map( A1 => n16280, A2 => n16243, ZN => n13889);
   U506 : INV_X4 port map( A => n13815, ZN => n13895);
   U507 : NAND2_X4 port map( A1 => n16289, A2 => n16285, ZN => n13815);
   U508 : INV_X4 port map( A => n13821, ZN => n13898);
   U509 : NAND2_X4 port map( A1 => n16286, A2 => n16285, ZN => n13821);
   U510 : INV_X4 port map( A => n13893, ZN => n13813);
   U511 : NAND2_X4 port map( A1 => n16285, A2 => n16290, ZN => n13893);
   U512 : INV_X4 port map( A => n13896, ZN => n13819);
   U513 : NAND2_X4 port map( A1 => n16283, A2 => n16285, ZN => n13896);
   U514 : INV_X4 port map( A => n11867, ZN => n301);
   U515 : INV_X4 port map( A => n13809, ZN => n13892);
   U516 : NAND2_X4 port map( A1 => n16285, A2 => n16264, ZN => n13809);
   U517 : INV_X8 port map( A => n11866, ZN => n302);
   U518 : AND2_X4 port map( A1 => n16441, A2 => N3583, ZN => r3013_A_3_port);
   U519 : AND2_X4 port map( A1 => n16454, A2 => N3570, ZN => r3007_A_3_port);
   U520 : AND2_X1 port map( A1 => n16285, A2 => n16243, ZN => n13816);
   U521 : INV_X4 port map( A => n13816, ZN => n303);
   U522 : AND2_X1 port map( A1 => n16280, A2 => n16286, ZN => n13822);
   U523 : INV_X4 port map( A => n13822, ZN => n304);
   U524 : INV_X2 port map( A => n303, ZN => n13865);
   U525 : INV_X2 port map( A => n304, ZN => n13868);
   U526 : AND2_X4 port map( A1 => n16264, A2 => n16244, ZN => n13826);
   U527 : AND2_X4 port map( A1 => n16280, A2 => n16245, ZN => n13808);
   U528 : NAND2_X2 port map( A1 => n16058, A2 => n16059, ZN => n5163);
   U529 : NAND2_X2 port map( A1 => n15830, A2 => n15831, ZN => n5133);
   U530 : NAND2_X2 port map( A1 => n15602, A2 => n15603, ZN => n5103);
   U531 : NAND2_X2 port map( A1 => n15374, A2 => n15375, ZN => n5073);
   U532 : NAND2_X2 port map( A1 => n15146, A2 => n15147, ZN => n5043);
   U533 : NAND2_X2 port map( A1 => n14918, A2 => n14919, ZN => n5013);
   U534 : NAND2_X2 port map( A1 => n14690, A2 => n14691, ZN => n4983);
   U535 : NAND2_X2 port map( A1 => n14462, A2 => n14463, ZN => n4953);
   U536 : NAND2_X2 port map( A1 => n14234, A2 => n14235, ZN => n4923);
   U537 : NAND2_X2 port map( A1 => n14006, A2 => n14007, ZN => n4893);
   U538 : NAND2_X2 port map( A1 => n15906, A2 => n15907, ZN => n5143);
   U539 : NAND2_X2 port map( A1 => n15678, A2 => n15679, ZN => n5113);
   U540 : NAND2_X2 port map( A1 => n15450, A2 => n15451, ZN => n5083);
   U541 : NAND2_X2 port map( A1 => n15222, A2 => n15223, ZN => n5053);
   U542 : NAND2_X2 port map( A1 => n14994, A2 => n14995, ZN => n5023);
   U543 : NAND2_X2 port map( A1 => n14766, A2 => n14767, ZN => n4993);
   U544 : NAND2_X2 port map( A1 => n14538, A2 => n14539, ZN => n4963);
   U545 : NAND2_X2 port map( A1 => n14310, A2 => n14311, ZN => n4933);
   U546 : NAND2_X2 port map( A1 => n14082, A2 => n14083, ZN => n4903);
   U547 : NAND2_X2 port map( A1 => n13966, A2 => n13967, ZN => n4885);
   U548 : NAND2_X2 port map( A1 => n16254, A2 => n16255, ZN => n5196);
   U549 : NAND2_X2 port map( A1 => n15866, A2 => n15867, ZN => n5135);
   U550 : NAND2_X2 port map( A1 => n15638, A2 => n15639, ZN => n5105);
   U551 : NAND2_X2 port map( A1 => n15410, A2 => n15411, ZN => n5075);
   U552 : NAND2_X2 port map( A1 => n15182, A2 => n15183, ZN => n5045);
   U553 : NAND2_X2 port map( A1 => n14954, A2 => n14955, ZN => n5015);
   U554 : NAND2_X2 port map( A1 => n14726, A2 => n14727, ZN => n4985);
   U555 : NAND2_X2 port map( A1 => n14498, A2 => n14499, ZN => n4955);
   U556 : NAND2_X2 port map( A1 => n14270, A2 => n14271, ZN => n4925);
   U557 : NAND2_X2 port map( A1 => n14042, A2 => n14043, ZN => n4895);
   U558 : NAND2_X2 port map( A1 => n13930, A2 => n13931, ZN => n4883);
   U559 : NAND2_X2 port map( A1 => n16214, A2 => n16215, ZN => n5192);
   U560 : NAND2_X2 port map( A1 => n13882, A2 => n13883, ZN => n4875);
   U561 : NAND2_X2 port map( A1 => n16152, A2 => n16153, ZN => n5172);
   U562 : NAND2_X2 port map( A1 => n16000, A2 => n16001, ZN => n5152);
   U563 : NAND2_X2 port map( A1 => n15772, A2 => n15773, ZN => n5122);
   U564 : NAND2_X2 port map( A1 => n15544, A2 => n15545, ZN => n5092);
   U565 : NAND2_X2 port map( A1 => n15316, A2 => n15317, ZN => n5062);
   U566 : NAND2_X2 port map( A1 => n15088, A2 => n15089, ZN => n5032);
   U567 : NAND2_X2 port map( A1 => n14860, A2 => n14861, ZN => n5002);
   U568 : NAND2_X2 port map( A1 => n14632, A2 => n14633, ZN => n4972);
   U569 : NAND2_X2 port map( A1 => n14404, A2 => n14405, ZN => n4942);
   U570 : NAND2_X2 port map( A1 => n14176, A2 => n14177, ZN => n4912);
   U571 : NAND2_X2 port map( A1 => n13797, A2 => n13798, ZN => n4871);
   U572 : NAND2_X2 port map( A1 => n16076, A2 => n16077, ZN => n5162);
   U573 : NAND2_X2 port map( A1 => n15924, A2 => n15925, ZN => n5142);
   U574 : NAND2_X2 port map( A1 => n15696, A2 => n15697, ZN => n5112);
   U575 : NAND2_X2 port map( A1 => n15468, A2 => n15469, ZN => n5082);
   U576 : NAND2_X2 port map( A1 => n15240, A2 => n15241, ZN => n5052);
   U577 : NAND2_X2 port map( A1 => n15012, A2 => n15013, ZN => n5022);
   U578 : NAND2_X2 port map( A1 => n14784, A2 => n14785, ZN => n4992);
   U579 : NAND2_X2 port map( A1 => n14556, A2 => n14557, ZN => n4962);
   U580 : NAND2_X2 port map( A1 => n14328, A2 => n14329, ZN => n4932);
   U581 : NAND2_X2 port map( A1 => n14100, A2 => n14101, ZN => n4902);
   U582 : NAND2_X2 port map( A1 => n15848, A2 => n15849, ZN => n5132);
   U583 : NAND2_X2 port map( A1 => n15620, A2 => n15621, ZN => n5102);
   U584 : NAND2_X2 port map( A1 => n15392, A2 => n15393, ZN => n5072);
   U585 : NAND2_X2 port map( A1 => n15164, A2 => n15165, ZN => n5042);
   U586 : NAND2_X2 port map( A1 => n14936, A2 => n14937, ZN => n5012);
   U587 : NAND2_X2 port map( A1 => n14708, A2 => n14709, ZN => n4982);
   U588 : NAND2_X2 port map( A1 => n14480, A2 => n14481, ZN => n4952);
   U589 : NAND2_X2 port map( A1 => n14252, A2 => n14253, ZN => n4922);
   U590 : NAND2_X2 port map( A1 => n14024, A2 => n14025, ZN => n4892);
   U591 : NAND2_X2 port map( A1 => n13948, A2 => n13949, ZN => n4882);
   U592 : NAND2_X2 port map( A1 => n16233, A2 => n16234, ZN => n5191);
   U593 : NAND2_X4 port map( A1 => n16287, A2 => n16281, ZN => n13810);
   U594 : NAND2_X4 port map( A1 => n16286, A2 => n16281, ZN => n13890);
   U595 : NOR3_X2 port map( A1 => CWP_4_port, A2 => CWP_5_port, A3 => 
                           CWP_3_port, ZN => n16281);
   U596 : NAND2_X2 port map( A1 => n13855_port, A2 => n13856_port, ZN => n4869)
                           ;
   U597 : NAND2_X2 port map( A1 => n16188, A2 => n16189, ZN => n5174);
   U598 : NAND2_X2 port map( A1 => n16036, A2 => n16037, ZN => n5154);
   U599 : NAND2_X2 port map( A1 => n15808, A2 => n15809, ZN => n5124);
   U600 : NAND2_X2 port map( A1 => n15580, A2 => n15581, ZN => n5094);
   U601 : NAND2_X2 port map( A1 => n15352, A2 => n15353, ZN => n5064);
   U602 : NAND2_X2 port map( A1 => n15124, A2 => n15125, ZN => n5034);
   U603 : NAND2_X2 port map( A1 => n14896, A2 => n14897, ZN => n5004);
   U604 : NAND2_X2 port map( A1 => n14668, A2 => n14669, ZN => n4974);
   U605 : NAND2_X2 port map( A1 => n14440, A2 => n14441, ZN => n4944);
   U606 : NAND2_X2 port map( A1 => n14212, A2 => n14213, ZN => n4914);
   U607 : AND2_X2 port map( A1 => n16245, A2 => n16244, ZN => n13871);
   U608 : AND2_X2 port map( A1 => n13630, A2 => n13629, ZN => n13498);
   U609 : AND2_X2 port map( A1 => n9919, A2 => n9917, ZN => n9788);
   U610 : AND2_X2 port map( A1 => n9035, A2 => n9032, ZN => n8903);
   U611 : AND2_X2 port map( A1 => n8146, A2 => n8143, ZN => n8014);
   U612 : AND4_X2 port map( A1 => n13780, A2 => n13628, A3 => n13331, A4 => 
                           n13781, ZN => n13647);
   U613 : INV_X2 port map( A => n16443, ZN => n16368);
   U614 : NAND3_X2 port map( A1 => n16433, A2 => WR, A3 => n16362, ZN => n16361
                           );
   U615 : INV_X4 port map( A => n13863, ZN => n13812);
   U616 : NAND2_X2 port map( A1 => n16264, A2 => n16281, ZN => n13863);
   U617 : AND2_X2 port map( A1 => n16441, A2 => N3584, ZN => r3013_A_4_port);
   U618 : AND2_X2 port map( A1 => N3572, A2 => n16454, ZN => ADD_RD1_5_port);
   U619 : NAND2_X2 port map( A1 => n16112, A2 => n16113, ZN => n5164);
   U620 : NAND2_X2 port map( A1 => n15960, A2 => n15961, ZN => n5144);
   U621 : NAND2_X2 port map( A1 => n15732, A2 => n15733, ZN => n5114);
   U622 : NAND2_X2 port map( A1 => n15504, A2 => n15505, ZN => n5084);
   U623 : NAND2_X2 port map( A1 => n15276, A2 => n15277, ZN => n5054);
   U624 : NAND2_X2 port map( A1 => n15048, A2 => n15049, ZN => n5024);
   U625 : NAND2_X2 port map( A1 => n14820, A2 => n14821, ZN => n4994);
   U626 : NAND2_X2 port map( A1 => n14592, A2 => n14593, ZN => n4964);
   U627 : NAND2_X2 port map( A1 => n14364, A2 => n14365, ZN => n4934);
   U628 : NAND2_X2 port map( A1 => n14136, A2 => n14137, ZN => n4904);
   U629 : NAND2_X2 port map( A1 => n13984, A2 => n13985, ZN => n4884);
   U630 : OAI22_X4 port map( A1 => n4800, A2 => n4809, B1 => n4839, B2 => n4808
                           , ZN => n4791);
   U631 : NOR3_X2 port map( A1 => n11865, A2 => n11866, A3 => n11864, ZN => 
                           n10226);
   U632 : INV_X2 port map( A => n4800, ZN => n4789);
   U633 : AND2_X2 port map( A1 => n16280, A2 => n16264, ZN => n13917);
   U634 : AND4_X2 port map( A1 => n13628, A2 => n13629, A3 => n11849, A4 => 
                           n13331, ZN => n13495);
   U635 : AND4_X2 port map( A1 => n9916, A2 => n9917, A3 => n9475, A4 => n9623,
                           ZN => n9783);
   U636 : AND4_X2 port map( A1 => n9031, A2 => n9032, A3 => n8586, A4 => n8735,
                           ZN => n8899);
   U637 : AND4_X2 port map( A1 => n8142, A2 => n8143, A3 => n7698, A4 => n7847,
                           ZN => n8010);
   U638 : NAND2_X2 port map( A1 => n5760, A2 => n5761, ZN => n5535);
   U639 : AND2_X2 port map( A1 => n5354, A2 => n5355, ZN => n5221);
   U640 : AND2_X2 port map( A1 => n5510, A2 => n5511, ZN => n5377);
   U641 : AND2_X2 port map( A1 => n7994, A2 => n7995, ZN => n7863);
   U642 : AND2_X2 port map( A1 => n7109, A2 => n7110, ZN => n6978);
   U643 : AND2_X2 port map( A1 => n6668, A2 => n6669, ZN => n6536);
   U644 : AND2_X2 port map( A1 => n6518, A2 => n6519, ZN => n6386);
   U645 : AND2_X2 port map( A1 => n6365, A2 => n6366, ZN => n6233);
   U646 : AND2_X2 port map( A1 => n6212, A2 => n6213, ZN => n6083);
   U647 : AND2_X2 port map( A1 => n6064, A2 => n6065, ZN => n5931);
   U648 : AND2_X2 port map( A1 => n5913, A2 => n5914, ZN => n5780);
   U649 : INV_X2 port map( A => n16430, ZN => n16364);
   U650 : NAND3_X2 port map( A1 => n16445, A2 => WR, A3 => n16366, ZN => n16365
                           );
   U651 : AND2_X2 port map( A1 => n13630, A2 => n13780, ZN => n13651);
   U652 : INV_X4 port map( A => n13869, ZN => n13824);
   U653 : NAND2_X2 port map( A1 => n16285, A2 => n16245, ZN => n13869);
   U654 : INV_X4 port map( A => n13866, ZN => n13818);
   U655 : NAND2_X2 port map( A1 => n16289, A2 => n16281, ZN => n13866);
   U656 : AND2_X2 port map( A1 => RD2, A2 => ENABLE, ZN => n16362);
   U657 : AND2_X2 port map( A1 => RD1, A2 => ENABLE, ZN => n16366);
   U658 : AND2_X2 port map( A1 => n16307, A2 => n16314, ZN => n13796);
   U659 : INV_X2 port map( A => ENABLE, ZN => n4786);
   U660 : AND2_X2 port map( A1 => n16454, A2 => N3571, ZN => r3007_A_4_port);
   U661 : AND2_X2 port map( A1 => N3585, A2 => n16441, ZN => ADD_RD2_5_port);
   U662 : INV_X2 port map( A => n5747, ZN => n5169);
   U663 : INV_X2 port map( A => n5740, ZN => n5159);
   U664 : INV_X2 port map( A => n5733, ZN => n5149);
   U665 : INV_X2 port map( A => n5726, ZN => n5139);
   U666 : INV_X2 port map( A => n5719, ZN => n5129);
   U667 : INV_X2 port map( A => n5712, ZN => n5119);
   U668 : INV_X2 port map( A => n5705, ZN => n5109);
   U669 : INV_X2 port map( A => n5698, ZN => n5099);
   U670 : INV_X2 port map( A => n5691, ZN => n5089);
   U671 : INV_X2 port map( A => n5684, ZN => n5079);
   U672 : INV_X2 port map( A => n5677, ZN => n5069);
   U673 : INV_X2 port map( A => n5670, ZN => n5059);
   U674 : INV_X2 port map( A => n5663, ZN => n5049);
   U675 : INV_X2 port map( A => n5656, ZN => n5039);
   U676 : INV_X2 port map( A => n5649, ZN => n5029);
   U677 : INV_X2 port map( A => n5642, ZN => n5019);
   U678 : INV_X2 port map( A => n5635, ZN => n5009);
   U679 : INV_X2 port map( A => n5628, ZN => n4999);
   U680 : INV_X2 port map( A => n5621, ZN => n4989);
   U681 : INV_X2 port map( A => n5614, ZN => n4979);
   U682 : INV_X2 port map( A => n5607, ZN => n4969);
   U683 : INV_X2 port map( A => n5600, ZN => n4959);
   U684 : INV_X2 port map( A => n5593, ZN => n4949);
   U685 : INV_X2 port map( A => n5586, ZN => n4939);
   U686 : INV_X2 port map( A => n5579, ZN => n4929);
   U687 : INV_X2 port map( A => n5572, ZN => n4919);
   U688 : INV_X2 port map( A => n5565, ZN => n4909);
   U689 : INV_X2 port map( A => n5558, ZN => n4899);
   U690 : INV_X2 port map( A => n5551, ZN => n4889);
   U691 : INV_X2 port map( A => n5544, ZN => n4879);
   U692 : INV_X2 port map( A => n5754, ZN => n5179);
   U693 : INV_X2 port map( A => n5536, ZN => n4863);
   U694 : INV_X2 port map( A => n5744, ZN => n5171);
   U695 : INV_X2 port map( A => n5737, ZN => n5161);
   U696 : INV_X2 port map( A => n5730, ZN => n5151);
   U697 : INV_X2 port map( A => n5723, ZN => n5141);
   U698 : INV_X2 port map( A => n5716, ZN => n5131);
   U699 : INV_X2 port map( A => n5709, ZN => n5121);
   U700 : INV_X2 port map( A => n5702, ZN => n5111);
   U701 : INV_X2 port map( A => n5695, ZN => n5101);
   U702 : INV_X2 port map( A => n5688, ZN => n5091);
   U703 : INV_X2 port map( A => n5681, ZN => n5081);
   U704 : INV_X2 port map( A => n5674, ZN => n5071);
   U705 : INV_X2 port map( A => n5667, ZN => n5061);
   U706 : INV_X2 port map( A => n5660, ZN => n5051);
   U707 : INV_X2 port map( A => n5653, ZN => n5041);
   U708 : INV_X2 port map( A => n5646, ZN => n5031);
   U709 : INV_X2 port map( A => n5639, ZN => n5021);
   U710 : INV_X2 port map( A => n5632, ZN => n5011);
   U711 : INV_X2 port map( A => n5625, ZN => n5001);
   U712 : INV_X2 port map( A => n5618, ZN => n4991);
   U713 : INV_X2 port map( A => n5611, ZN => n4981);
   U714 : INV_X2 port map( A => n5604, ZN => n4971);
   U715 : INV_X2 port map( A => n5597, ZN => n4961);
   U716 : INV_X2 port map( A => n5590, ZN => n4951);
   U717 : INV_X2 port map( A => n5583, ZN => n4941);
   U718 : INV_X2 port map( A => n5576, ZN => n4931);
   U719 : INV_X2 port map( A => n5569, ZN => n4921);
   U720 : INV_X2 port map( A => n5562, ZN => n4911);
   U721 : INV_X2 port map( A => n5555, ZN => n4901);
   U722 : INV_X2 port map( A => n5548, ZN => n4891);
   U723 : INV_X2 port map( A => n5541, ZN => n4881);
   U724 : INV_X2 port map( A => n5531, ZN => n4867);
   U725 : INV_X2 port map( A => n5751, ZN => n5181);
   U726 : NAND2_X2 port map( A1 => n15884, A2 => n15885, ZN => n5134);
   U727 : NAND2_X2 port map( A1 => n15656, A2 => n15657, ZN => n5104);
   U728 : NAND2_X2 port map( A1 => n15428, A2 => n15429, ZN => n5074);
   U729 : NAND2_X2 port map( A1 => n15200, A2 => n15201, ZN => n5044);
   U730 : NAND2_X2 port map( A1 => n14972, A2 => n14973, ZN => n5014);
   U731 : NAND2_X2 port map( A1 => n14744, A2 => n14745, ZN => n4984);
   U732 : NAND2_X2 port map( A1 => n14516, A2 => n14517, ZN => n4954);
   U733 : NAND2_X2 port map( A1 => n14288, A2 => n14289, ZN => n4924);
   U734 : NAND2_X2 port map( A1 => n14060, A2 => n14061, ZN => n4894);
   U735 : NAND2_X2 port map( A1 => n13907, A2 => n13908, ZN => n4873);
   U736 : NAND2_X2 port map( A1 => n16273, A2 => n16274, ZN => n5195);
   U737 : INV_X2 port map( A => RESET, ZN => n5368);
   U738 : OR3_X1 port map( A1 => n4802, A2 => n4811, A3 => n4839, ZN => n4792);
   U739 : INV_X2 port map( A => n4792, ZN => n305);
   U740 : BUF_X1 port map( A => CLK, Z => n1003);
   U741 : BUF_X1 port map( A => CLK, Z => n984);
   U742 : BUF_X1 port map( A => CLK, Z => n997);
   U743 : BUF_X1 port map( A => CLK, Z => n1002);
   U744 : BUF_X1 port map( A => CLK, Z => n1001);
   U745 : BUF_X1 port map( A => CLK, Z => n987);
   U746 : BUF_X1 port map( A => CLK, Z => n998);
   U747 : BUF_X1 port map( A => CLK, Z => n1000);
   U748 : BUF_X1 port map( A => CLK, Z => n999);
   U749 : BUF_X1 port map( A => CLK, Z => n985);
   U750 : BUF_X1 port map( A => CLK, Z => n995);
   U751 : BUF_X1 port map( A => CLK, Z => n994);
   U752 : BUF_X1 port map( A => CLK, Z => n993);
   U753 : BUF_X1 port map( A => CLK, Z => n992);
   U754 : BUF_X1 port map( A => CLK, Z => n991);
   U755 : BUF_X1 port map( A => CLK, Z => n988);
   U756 : BUF_X1 port map( A => CLK, Z => n990);
   U757 : BUF_X1 port map( A => CLK, Z => n989);
   U758 : BUF_X1 port map( A => CLK, Z => n996);
   U759 : BUF_X1 port map( A => CLK, Z => n986);
   U760 : BUF_X1 port map( A => CLK, Z => n983);
   U761 : BUF_X1 port map( A => CLK, Z => n982);
   U762 : BUF_X1 port map( A => r3007_A_1_port, Z => n723);
   U763 : BUF_X1 port map( A => r3007_A_1_port, Z => n724);
   U764 : BUF_X1 port map( A => r3007_A_1_port, Z => n725);
   U765 : BUF_X1 port map( A => r3007_A_1_port, Z => n726);
   U766 : BUF_X1 port map( A => r3007_A_1_port, Z => n727);
   U767 : BUF_X1 port map( A => r3007_A_1_port, Z => n728);
   U768 : BUF_X1 port map( A => r3007_A_1_port, Z => n729);
   U769 : BUF_X1 port map( A => r3007_A_1_port, Z => n730);
   U770 : BUF_X1 port map( A => r3013_A_1_port, Z => n637);
   U771 : BUF_X1 port map( A => r3013_A_1_port, Z => n638);
   U772 : BUF_X1 port map( A => r3013_A_1_port, Z => n639);
   U773 : BUF_X1 port map( A => r3013_A_1_port, Z => n640);
   U774 : BUF_X1 port map( A => r3013_A_1_port, Z => n641);
   U775 : BUF_X1 port map( A => r3013_A_1_port, Z => n642);
   U776 : BUF_X1 port map( A => r3013_A_1_port, Z => n643);
   U777 : BUF_X1 port map( A => r3013_A_1_port, Z => n644);
   U778 : BUF_X1 port map( A => r3007_A_1_port, Z => n731);
   U779 : BUF_X1 port map( A => r3013_A_1_port, Z => n645);
   U780 : BUF_X2 port map( A => SWP_4_port, Z => n841);
   U781 : BUF_X2 port map( A => SWP_5_port, Z => n846);
   U782 : BUF_X2 port map( A => SWP_4_port, Z => n844);
   U783 : BUF_X2 port map( A => SWP_5_port, Z => n848);
   U784 : BUF_X2 port map( A => SWP_4_port, Z => n843);
   U785 : BUF_X2 port map( A => SWP_4_port, Z => n842);
   U786 : BUF_X2 port map( A => SWP_5_port, Z => n847);
   U787 : BUF_X1 port map( A => SWP_5_port, Z => n849);
   U788 : BUF_X1 port map( A => SWP_4_port, Z => n845);
   U789 : XNOR2_X1 port map( A => WR_ADD(4), B => sub_65_carry_4_port, ZN => 
                           N3592);
   U790 : NAND2_X1 port map( A1 => n1004, A2 => N3590, ZN => 
                           sub_65_carry_4_port);
   U791 : INV_X1 port map( A => WR_ADD(3), ZN => n1004);
   U792 : XNOR2_X1 port map( A => RD1_ADD(4), B => sub_63_carry_4_port, ZN => 
                           N3566);
   U793 : NAND2_X1 port map( A1 => n1006, A2 => N3564, ZN => 
                           sub_63_carry_4_port);
   U794 : INV_X1 port map( A => RD1_ADD(3), ZN => n1006);
   U795 : XNOR2_X1 port map( A => RD2_ADD(4), B => sub_64_carry_4_port, ZN => 
                           N3579);
   U796 : NAND2_X1 port map( A1 => n1005, A2 => N3577, ZN => 
                           sub_64_carry_4_port);
   U797 : INV_X1 port map( A => RD2_ADD(3), ZN => n1005);
   U798 : XNOR2_X1 port map( A => WR_ADD(3), B => WR_ADD(2), ZN => N3591);
   U799 : XNOR2_X1 port map( A => RD1_ADD(3), B => RD1_ADD(2), ZN => N3565);
   U800 : XNOR2_X1 port map( A => RD2_ADD(3), B => RD2_ADD(2), ZN => N3578);
   U801 : BUF_X1 port map( A => SWP_0_port, Z => n807);
   U802 : BUF_X1 port map( A => SWP_0_port, Z => n808);
   U803 : BUF_X1 port map( A => SWP_0_port, Z => n805);
   U804 : BUF_X1 port map( A => SWP_0_port, Z => n806);
   U805 : BUF_X1 port map( A => SWP_0_port, Z => n812);
   U806 : BUF_X1 port map( A => SWP_0_port, Z => n809);
   U807 : BUF_X1 port map( A => SWP_0_port, Z => n810);
   U808 : BUF_X1 port map( A => SWP_0_port, Z => n811);
   U809 : BUF_X1 port map( A => SWP_0_port, Z => n813);
   U810 : CLKBUF_X1 port map( A => n13803, Z => n306);
   U811 : CLKBUF_X1 port map( A => n13803, Z => n307);
   U812 : CLKBUF_X1 port map( A => n13803, Z => n308);
   U813 : CLKBUF_X1 port map( A => n13803, Z => n309);
   U814 : CLKBUF_X1 port map( A => n13803, Z => n310);
   U815 : CLKBUF_X1 port map( A => n13803, Z => n311);
   U816 : CLKBUF_X1 port map( A => n13803, Z => n312);
   U817 : CLKBUF_X1 port map( A => n13803, Z => n313);
   U818 : CLKBUF_X1 port map( A => n13803, Z => n314);
   U819 : CLKBUF_X1 port map( A => n13803, Z => n315);
   U820 : CLKBUF_X1 port map( A => n13803, Z => n316);
   U821 : CLKBUF_X1 port map( A => n13804, Z => n317);
   U822 : CLKBUF_X1 port map( A => n13804, Z => n318);
   U823 : CLKBUF_X1 port map( A => n13804, Z => n319);
   U824 : CLKBUF_X1 port map( A => n13804, Z => n320);
   U825 : CLKBUF_X1 port map( A => n13804, Z => n321);
   U826 : CLKBUF_X1 port map( A => n13804, Z => n322);
   U827 : CLKBUF_X1 port map( A => n13804, Z => n323);
   U828 : CLKBUF_X1 port map( A => n13804, Z => n324);
   U829 : CLKBUF_X1 port map( A => n13804, Z => n325);
   U830 : CLKBUF_X1 port map( A => n13804, Z => n326);
   U831 : CLKBUF_X1 port map( A => n13804, Z => n327);
   U832 : CLKBUF_X1 port map( A => n13806, Z => n328);
   U833 : CLKBUF_X1 port map( A => n13806, Z => n329);
   U834 : CLKBUF_X1 port map( A => n13806, Z => n330);
   U835 : CLKBUF_X1 port map( A => n13806, Z => n331);
   U836 : CLKBUF_X1 port map( A => n13806, Z => n332);
   U837 : CLKBUF_X1 port map( A => n13806, Z => n333);
   U838 : CLKBUF_X1 port map( A => n13806, Z => n334);
   U839 : CLKBUF_X1 port map( A => n13806, Z => n335);
   U840 : CLKBUF_X1 port map( A => n13806, Z => n336);
   U841 : CLKBUF_X1 port map( A => n13806, Z => n337);
   U842 : CLKBUF_X1 port map( A => n13806, Z => n338);
   U843 : CLKBUF_X1 port map( A => n13814, Z => n339);
   U844 : CLKBUF_X1 port map( A => n13814, Z => n340);
   U845 : CLKBUF_X1 port map( A => n13814, Z => n341);
   U846 : CLKBUF_X1 port map( A => n13814, Z => n342);
   U847 : CLKBUF_X1 port map( A => n13814, Z => n343);
   U848 : CLKBUF_X1 port map( A => n13814, Z => n344);
   U849 : CLKBUF_X1 port map( A => n13814, Z => n345);
   U850 : CLKBUF_X1 port map( A => n13814, Z => n346);
   U851 : CLKBUF_X1 port map( A => n13814, Z => n347);
   U852 : CLKBUF_X1 port map( A => n13814, Z => n348);
   U853 : CLKBUF_X1 port map( A => n13814, Z => n349);
   U854 : CLKBUF_X1 port map( A => n13820, Z => n350);
   U855 : CLKBUF_X1 port map( A => n13820, Z => n351);
   U856 : CLKBUF_X1 port map( A => n13820, Z => n352);
   U857 : CLKBUF_X1 port map( A => n13820, Z => n353);
   U858 : CLKBUF_X1 port map( A => n13820, Z => n354);
   U859 : CLKBUF_X1 port map( A => n13820, Z => n355);
   U860 : CLKBUF_X1 port map( A => n13820, Z => n356);
   U861 : CLKBUF_X1 port map( A => n13820, Z => n357);
   U862 : CLKBUF_X1 port map( A => n13820, Z => n358);
   U863 : CLKBUF_X1 port map( A => n13820, Z => n359);
   U864 : CLKBUF_X1 port map( A => n13820, Z => n360);
   U865 : CLKBUF_X1 port map( A => n13831_port, Z => n361);
   U866 : CLKBUF_X1 port map( A => n13831_port, Z => n362);
   U867 : CLKBUF_X1 port map( A => n13831_port, Z => n363);
   U868 : CLKBUF_X1 port map( A => n13831_port, Z => n364);
   U869 : CLKBUF_X1 port map( A => n13831_port, Z => n365);
   U870 : CLKBUF_X1 port map( A => n13831_port, Z => n366);
   U871 : CLKBUF_X1 port map( A => n13831_port, Z => n367);
   U872 : CLKBUF_X1 port map( A => n13831_port, Z => n368);
   U873 : CLKBUF_X1 port map( A => n13831_port, Z => n369);
   U874 : CLKBUF_X1 port map( A => n13831_port, Z => n370);
   U875 : CLKBUF_X1 port map( A => n13831_port, Z => n371);
   U876 : CLKBUF_X1 port map( A => n13832_port, Z => n372);
   U877 : CLKBUF_X1 port map( A => n13832_port, Z => n373);
   U878 : CLKBUF_X1 port map( A => n13832_port, Z => n374);
   U879 : CLKBUF_X1 port map( A => n13832_port, Z => n375);
   U880 : CLKBUF_X1 port map( A => n13832_port, Z => n376);
   U881 : CLKBUF_X1 port map( A => n13832_port, Z => n377);
   U882 : CLKBUF_X1 port map( A => n13832_port, Z => n378);
   U883 : CLKBUF_X1 port map( A => n13832_port, Z => n379);
   U884 : CLKBUF_X1 port map( A => n13832_port, Z => n380);
   U885 : CLKBUF_X1 port map( A => n13832_port, Z => n381);
   U886 : CLKBUF_X1 port map( A => n13832_port, Z => n382);
   U887 : CLKBUF_X1 port map( A => n13834_port, Z => n383);
   U888 : CLKBUF_X1 port map( A => n13834_port, Z => n384);
   U889 : CLKBUF_X1 port map( A => n13834_port, Z => n385);
   U890 : CLKBUF_X1 port map( A => n13834_port, Z => n386);
   U891 : CLKBUF_X1 port map( A => n13834_port, Z => n387);
   U892 : CLKBUF_X1 port map( A => n13834_port, Z => n388);
   U893 : CLKBUF_X1 port map( A => n13834_port, Z => n389);
   U894 : CLKBUF_X1 port map( A => n13834_port, Z => n390);
   U895 : CLKBUF_X1 port map( A => n13834_port, Z => n391);
   U896 : CLKBUF_X1 port map( A => n13834_port, Z => n392);
   U897 : CLKBUF_X1 port map( A => n13834_port, Z => n393);
   U898 : CLKBUF_X1 port map( A => n13835_port, Z => n394);
   U899 : CLKBUF_X1 port map( A => n13835_port, Z => n395);
   U900 : CLKBUF_X1 port map( A => n13835_port, Z => n396);
   U901 : CLKBUF_X1 port map( A => n13835_port, Z => n397);
   U902 : CLKBUF_X1 port map( A => n13835_port, Z => n398);
   U903 : CLKBUF_X1 port map( A => n13835_port, Z => n399);
   U904 : CLKBUF_X1 port map( A => n13835_port, Z => n400);
   U905 : CLKBUF_X1 port map( A => n13835_port, Z => n401);
   U906 : CLKBUF_X1 port map( A => n13835_port, Z => n402);
   U907 : CLKBUF_X1 port map( A => n13835_port, Z => n403);
   U908 : CLKBUF_X1 port map( A => n13835_port, Z => n404);
   U909 : CLKBUF_X1 port map( A => n13836_port, Z => n405);
   U910 : CLKBUF_X1 port map( A => n13836_port, Z => n406);
   U911 : CLKBUF_X1 port map( A => n13836_port, Z => n407);
   U912 : CLKBUF_X1 port map( A => n13836_port, Z => n408);
   U913 : CLKBUF_X1 port map( A => n13836_port, Z => n409);
   U914 : CLKBUF_X1 port map( A => n13836_port, Z => n410);
   U915 : CLKBUF_X1 port map( A => n13836_port, Z => n411);
   U916 : CLKBUF_X1 port map( A => n13836_port, Z => n412);
   U917 : CLKBUF_X1 port map( A => n13836_port, Z => n413);
   U918 : CLKBUF_X1 port map( A => n13836_port, Z => n414);
   U919 : CLKBUF_X1 port map( A => n13836_port, Z => n415);
   U920 : CLKBUF_X1 port map( A => n13837_port, Z => n416);
   U921 : CLKBUF_X1 port map( A => n13837_port, Z => n417);
   U922 : CLKBUF_X1 port map( A => n13837_port, Z => n418);
   U923 : CLKBUF_X1 port map( A => n13837_port, Z => n419);
   U924 : CLKBUF_X1 port map( A => n13837_port, Z => n420);
   U925 : CLKBUF_X1 port map( A => n13837_port, Z => n421);
   U926 : CLKBUF_X1 port map( A => n13837_port, Z => n422);
   U927 : CLKBUF_X1 port map( A => n13837_port, Z => n423);
   U928 : CLKBUF_X1 port map( A => n13837_port, Z => n424);
   U929 : CLKBUF_X1 port map( A => n13837_port, Z => n425);
   U930 : CLKBUF_X1 port map( A => n13837_port, Z => n426);
   U931 : CLKBUF_X1 port map( A => n13838_port, Z => n427);
   U932 : CLKBUF_X1 port map( A => n13838_port, Z => n428);
   U933 : CLKBUF_X1 port map( A => n13838_port, Z => n429);
   U934 : CLKBUF_X1 port map( A => n13838_port, Z => n430);
   U935 : CLKBUF_X1 port map( A => n13838_port, Z => n431);
   U936 : CLKBUF_X1 port map( A => n13838_port, Z => n432);
   U937 : CLKBUF_X1 port map( A => n13838_port, Z => n433);
   U938 : CLKBUF_X1 port map( A => n13838_port, Z => n434);
   U939 : CLKBUF_X1 port map( A => n13838_port, Z => n435);
   U940 : CLKBUF_X1 port map( A => n13838_port, Z => n436);
   U941 : CLKBUF_X1 port map( A => n13838_port, Z => n437);
   U942 : CLKBUF_X1 port map( A => n13840_port, Z => n438);
   U943 : CLKBUF_X1 port map( A => n13840_port, Z => n439);
   U944 : CLKBUF_X1 port map( A => n13840_port, Z => n440);
   U945 : CLKBUF_X1 port map( A => n13840_port, Z => n441);
   U946 : CLKBUF_X1 port map( A => n13840_port, Z => n442);
   U947 : CLKBUF_X1 port map( A => n13840_port, Z => n443);
   U948 : CLKBUF_X1 port map( A => n13840_port, Z => n444);
   U949 : CLKBUF_X1 port map( A => n13840_port, Z => n445);
   U950 : CLKBUF_X1 port map( A => n13840_port, Z => n446);
   U951 : CLKBUF_X1 port map( A => n13840_port, Z => n447);
   U952 : CLKBUF_X1 port map( A => n13840_port, Z => n448);
   U953 : CLKBUF_X1 port map( A => n13841_port, Z => n449);
   U954 : CLKBUF_X1 port map( A => n13841_port, Z => n450);
   U955 : CLKBUF_X1 port map( A => n13841_port, Z => n451);
   U956 : CLKBUF_X1 port map( A => n13841_port, Z => n452);
   U957 : CLKBUF_X1 port map( A => n13841_port, Z => n453);
   U958 : CLKBUF_X1 port map( A => n13841_port, Z => n454);
   U959 : CLKBUF_X1 port map( A => n13841_port, Z => n455);
   U960 : CLKBUF_X1 port map( A => n13841_port, Z => n456);
   U961 : CLKBUF_X1 port map( A => n13841_port, Z => n457);
   U962 : CLKBUF_X1 port map( A => n13841_port, Z => n458);
   U963 : CLKBUF_X1 port map( A => n13841_port, Z => n459);
   U964 : CLKBUF_X1 port map( A => n13842_port, Z => n460);
   U965 : CLKBUF_X1 port map( A => n13842_port, Z => n461);
   U966 : CLKBUF_X1 port map( A => n13842_port, Z => n462);
   U967 : CLKBUF_X1 port map( A => n13842_port, Z => n463);
   U968 : CLKBUF_X1 port map( A => n13842_port, Z => n464);
   U969 : CLKBUF_X1 port map( A => n13842_port, Z => n465);
   U970 : CLKBUF_X1 port map( A => n13842_port, Z => n466);
   U971 : CLKBUF_X1 port map( A => n13842_port, Z => n467);
   U972 : CLKBUF_X1 port map( A => n13842_port, Z => n468);
   U973 : CLKBUF_X1 port map( A => n13842_port, Z => n469);
   U974 : CLKBUF_X1 port map( A => n13842_port, Z => n470);
   U975 : CLKBUF_X1 port map( A => n13843_port, Z => n471);
   U976 : CLKBUF_X1 port map( A => n13843_port, Z => n472);
   U977 : CLKBUF_X1 port map( A => n13843_port, Z => n473);
   U978 : CLKBUF_X1 port map( A => n13843_port, Z => n474);
   U979 : CLKBUF_X1 port map( A => n13843_port, Z => n475);
   U980 : CLKBUF_X1 port map( A => n13843_port, Z => n476);
   U981 : CLKBUF_X1 port map( A => n13843_port, Z => n477);
   U982 : CLKBUF_X1 port map( A => n13843_port, Z => n478);
   U983 : CLKBUF_X1 port map( A => n13843_port, Z => n479);
   U984 : CLKBUF_X1 port map( A => n13843_port, Z => n480);
   U985 : CLKBUF_X1 port map( A => n13843_port, Z => n481);
   U986 : CLKBUF_X1 port map( A => n13844_port, Z => n482);
   U987 : CLKBUF_X1 port map( A => n13844_port, Z => n483);
   U988 : CLKBUF_X1 port map( A => n13844_port, Z => n484);
   U989 : CLKBUF_X1 port map( A => n13844_port, Z => n485);
   U990 : CLKBUF_X1 port map( A => n13844_port, Z => n486);
   U991 : CLKBUF_X1 port map( A => n13844_port, Z => n487);
   U992 : CLKBUF_X1 port map( A => n13844_port, Z => n488);
   U993 : CLKBUF_X1 port map( A => n13844_port, Z => n489);
   U994 : CLKBUF_X1 port map( A => n13844_port, Z => n490);
   U995 : CLKBUF_X1 port map( A => n13844_port, Z => n491);
   U996 : CLKBUF_X1 port map( A => n13844_port, Z => n492);
   U997 : CLKBUF_X1 port map( A => n13846_port, Z => n493);
   U998 : CLKBUF_X1 port map( A => n13846_port, Z => n494);
   U999 : CLKBUF_X1 port map( A => n13846_port, Z => n495);
   U1000 : CLKBUF_X1 port map( A => n13846_port, Z => n496);
   U1001 : CLKBUF_X1 port map( A => n13846_port, Z => n497);
   U1002 : CLKBUF_X1 port map( A => n13846_port, Z => n498);
   U1003 : CLKBUF_X1 port map( A => n13846_port, Z => n499);
   U1004 : CLKBUF_X1 port map( A => n13846_port, Z => n500);
   U1005 : CLKBUF_X1 port map( A => n13846_port, Z => n501);
   U1006 : CLKBUF_X1 port map( A => n13846_port, Z => n502);
   U1007 : CLKBUF_X1 port map( A => n13846_port, Z => n503);
   U1008 : CLKBUF_X1 port map( A => n13847_port, Z => n504);
   U1009 : CLKBUF_X1 port map( A => n13847_port, Z => n505);
   U1010 : CLKBUF_X1 port map( A => n13847_port, Z => n506);
   U1011 : CLKBUF_X1 port map( A => n13847_port, Z => n507);
   U1012 : CLKBUF_X1 port map( A => n13847_port, Z => n508);
   U1013 : CLKBUF_X1 port map( A => n13847_port, Z => n509);
   U1014 : CLKBUF_X1 port map( A => n13847_port, Z => n510);
   U1015 : CLKBUF_X1 port map( A => n13847_port, Z => n511);
   U1016 : CLKBUF_X1 port map( A => n13847_port, Z => n512);
   U1017 : CLKBUF_X1 port map( A => n13847_port, Z => n513);
   U1018 : CLKBUF_X1 port map( A => n13847_port, Z => n514);
   U1019 : CLKBUF_X1 port map( A => n13848_port, Z => n515);
   U1020 : CLKBUF_X1 port map( A => n13848_port, Z => n516);
   U1021 : CLKBUF_X1 port map( A => n13848_port, Z => n517);
   U1022 : CLKBUF_X1 port map( A => n13848_port, Z => n518);
   U1023 : CLKBUF_X1 port map( A => n13848_port, Z => n519);
   U1024 : CLKBUF_X1 port map( A => n13848_port, Z => n520);
   U1025 : CLKBUF_X1 port map( A => n13848_port, Z => n521);
   U1026 : CLKBUF_X1 port map( A => n13848_port, Z => n522);
   U1027 : CLKBUF_X1 port map( A => n13848_port, Z => n523);
   U1028 : CLKBUF_X1 port map( A => n13848_port, Z => n524);
   U1029 : CLKBUF_X1 port map( A => n13848_port, Z => n525);
   U1030 : CLKBUF_X1 port map( A => n13849_port, Z => n526);
   U1031 : CLKBUF_X1 port map( A => n13849_port, Z => n527);
   U1032 : CLKBUF_X1 port map( A => n13849_port, Z => n528);
   U1033 : CLKBUF_X1 port map( A => n13849_port, Z => n529);
   U1034 : CLKBUF_X1 port map( A => n13849_port, Z => n530);
   U1035 : CLKBUF_X1 port map( A => n13849_port, Z => n531);
   U1036 : CLKBUF_X1 port map( A => n13849_port, Z => n532);
   U1037 : CLKBUF_X1 port map( A => n13849_port, Z => n533);
   U1038 : CLKBUF_X1 port map( A => n13849_port, Z => n534);
   U1039 : CLKBUF_X1 port map( A => n13849_port, Z => n535);
   U1040 : CLKBUF_X1 port map( A => n13849_port, Z => n536);
   U1041 : CLKBUF_X1 port map( A => n13850_port, Z => n537);
   U1042 : CLKBUF_X1 port map( A => n13850_port, Z => n538);
   U1043 : CLKBUF_X1 port map( A => n13850_port, Z => n539);
   U1044 : CLKBUF_X1 port map( A => n13850_port, Z => n540);
   U1045 : CLKBUF_X1 port map( A => n13850_port, Z => n541);
   U1046 : CLKBUF_X1 port map( A => n13850_port, Z => n542);
   U1047 : CLKBUF_X1 port map( A => n13850_port, Z => n543);
   U1048 : CLKBUF_X1 port map( A => n13850_port, Z => n544);
   U1049 : CLKBUF_X1 port map( A => n13850_port, Z => n545);
   U1050 : CLKBUF_X1 port map( A => n13850_port, Z => n546);
   U1051 : CLKBUF_X1 port map( A => n13850_port, Z => n547);
   U1052 : CLKBUF_X1 port map( A => n13852_port, Z => n548);
   U1053 : CLKBUF_X1 port map( A => n13852_port, Z => n549);
   U1054 : CLKBUF_X1 port map( A => n13852_port, Z => n550);
   U1055 : CLKBUF_X1 port map( A => n13852_port, Z => n551);
   U1056 : CLKBUF_X1 port map( A => n13852_port, Z => n552);
   U1057 : CLKBUF_X1 port map( A => n13852_port, Z => n553);
   U1058 : CLKBUF_X1 port map( A => n13852_port, Z => n554);
   U1059 : CLKBUF_X1 port map( A => n13852_port, Z => n555);
   U1060 : CLKBUF_X1 port map( A => n13852_port, Z => n556);
   U1061 : CLKBUF_X1 port map( A => n13852_port, Z => n557);
   U1062 : CLKBUF_X1 port map( A => n13852_port, Z => n558);
   U1063 : CLKBUF_X1 port map( A => n13853_port, Z => n559);
   U1064 : CLKBUF_X1 port map( A => n13853_port, Z => n560);
   U1065 : CLKBUF_X1 port map( A => n13853_port, Z => n561);
   U1066 : CLKBUF_X1 port map( A => n13853_port, Z => n562);
   U1067 : CLKBUF_X1 port map( A => n13853_port, Z => n563);
   U1068 : CLKBUF_X1 port map( A => n13853_port, Z => n564);
   U1069 : CLKBUF_X1 port map( A => n13853_port, Z => n565);
   U1070 : CLKBUF_X1 port map( A => n13853_port, Z => n566);
   U1071 : CLKBUF_X1 port map( A => n13853_port, Z => n567);
   U1072 : CLKBUF_X1 port map( A => n13853_port, Z => n568);
   U1073 : CLKBUF_X1 port map( A => n13853_port, Z => n569);
   U1074 : CLKBUF_X1 port map( A => n13854_port, Z => n570);
   U1075 : CLKBUF_X1 port map( A => n13854_port, Z => n571);
   U1076 : CLKBUF_X1 port map( A => n13854_port, Z => n572);
   U1077 : CLKBUF_X1 port map( A => n13854_port, Z => n573);
   U1078 : CLKBUF_X1 port map( A => n13854_port, Z => n574);
   U1079 : CLKBUF_X1 port map( A => n13854_port, Z => n575);
   U1080 : CLKBUF_X1 port map( A => n13854_port, Z => n576);
   U1081 : CLKBUF_X1 port map( A => n13854_port, Z => n577);
   U1082 : CLKBUF_X1 port map( A => n13854_port, Z => n578);
   U1083 : CLKBUF_X1 port map( A => n13854_port, Z => n579);
   U1084 : CLKBUF_X1 port map( A => n13854_port, Z => n580);
   U1085 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n581);
   U1086 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n582);
   U1087 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n583);
   U1088 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n584);
   U1089 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n585);
   U1090 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n586);
   U1091 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n587);
   U1092 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n588);
   U1093 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n589);
   U1094 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n590);
   U1095 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n591);
   U1096 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n592);
   U1097 : CLKBUF_X1 port map( A => r3013_A_2_port, Z => n593);
   U1098 : CLKBUF_X1 port map( A => n645, Z => n594);
   U1099 : CLKBUF_X1 port map( A => n645, Z => n595);
   U1100 : CLKBUF_X1 port map( A => n645, Z => n596);
   U1101 : CLKBUF_X1 port map( A => n644, Z => n597);
   U1102 : CLKBUF_X1 port map( A => n644, Z => n598);
   U1103 : CLKBUF_X1 port map( A => n644, Z => n599);
   U1104 : CLKBUF_X1 port map( A => n644, Z => n600);
   U1105 : CLKBUF_X1 port map( A => n644, Z => n601);
   U1106 : CLKBUF_X1 port map( A => n643, Z => n602);
   U1107 : CLKBUF_X1 port map( A => n643, Z => n603);
   U1108 : CLKBUF_X1 port map( A => n643, Z => n604);
   U1109 : CLKBUF_X1 port map( A => n643, Z => n605);
   U1110 : CLKBUF_X1 port map( A => n643, Z => n606);
   U1111 : CLKBUF_X1 port map( A => n642, Z => n607);
   U1112 : CLKBUF_X1 port map( A => n642, Z => n608);
   U1113 : CLKBUF_X1 port map( A => n642, Z => n609);
   U1114 : CLKBUF_X1 port map( A => n642, Z => n610);
   U1115 : CLKBUF_X1 port map( A => n642, Z => n611);
   U1116 : CLKBUF_X1 port map( A => n641, Z => n612);
   U1117 : CLKBUF_X1 port map( A => n641, Z => n613);
   U1118 : CLKBUF_X1 port map( A => n641, Z => n614);
   U1119 : CLKBUF_X1 port map( A => n641, Z => n615);
   U1120 : CLKBUF_X1 port map( A => n641, Z => n616);
   U1121 : CLKBUF_X1 port map( A => n640, Z => n617);
   U1122 : CLKBUF_X1 port map( A => n640, Z => n618);
   U1123 : CLKBUF_X1 port map( A => n640, Z => n619);
   U1124 : CLKBUF_X1 port map( A => n640, Z => n620);
   U1125 : CLKBUF_X1 port map( A => n640, Z => n621);
   U1126 : CLKBUF_X1 port map( A => n639, Z => n622);
   U1127 : CLKBUF_X1 port map( A => n639, Z => n623);
   U1128 : CLKBUF_X1 port map( A => n639, Z => n624);
   U1129 : CLKBUF_X1 port map( A => n639, Z => n625);
   U1130 : CLKBUF_X1 port map( A => n639, Z => n626);
   U1131 : CLKBUF_X1 port map( A => n638, Z => n627);
   U1132 : CLKBUF_X1 port map( A => n638, Z => n628);
   U1133 : CLKBUF_X1 port map( A => n638, Z => n629);
   U1134 : CLKBUF_X1 port map( A => n638, Z => n630);
   U1135 : CLKBUF_X1 port map( A => n638, Z => n631);
   U1136 : CLKBUF_X1 port map( A => n637, Z => n632);
   U1137 : CLKBUF_X1 port map( A => n637, Z => n633);
   U1138 : CLKBUF_X1 port map( A => n637, Z => n634);
   U1139 : CLKBUF_X1 port map( A => n637, Z => n635);
   U1140 : CLKBUF_X1 port map( A => n637, Z => n636);
   U1141 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n646);
   U1142 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n647);
   U1143 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n648);
   U1144 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n649);
   U1145 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n650);
   U1146 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n651);
   U1147 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n652);
   U1148 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n653);
   U1149 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n654);
   U1150 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n655);
   U1151 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n656);
   U1152 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n657);
   U1153 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n658);
   U1154 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n659);
   U1155 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n660);
   U1156 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n661);
   U1157 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n662);
   U1158 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n663);
   U1159 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n664);
   U1160 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n665);
   U1161 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n666);
   U1162 : CLKBUF_X1 port map( A => r3013_A_0_port, Z => n667);
   U1163 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n668);
   U1164 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n669);
   U1165 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n670);
   U1166 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n671);
   U1167 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n672);
   U1168 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n673);
   U1169 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n674);
   U1170 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n675);
   U1171 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n676);
   U1172 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n677);
   U1173 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n678);
   U1174 : CLKBUF_X1 port map( A => r3007_A_2_port, Z => n679);
   U1175 : CLKBUF_X1 port map( A => n731, Z => n680);
   U1176 : CLKBUF_X1 port map( A => n731, Z => n681);
   U1177 : CLKBUF_X1 port map( A => n731, Z => n682);
   U1178 : CLKBUF_X1 port map( A => n730, Z => n683);
   U1179 : CLKBUF_X1 port map( A => n730, Z => n684);
   U1180 : CLKBUF_X1 port map( A => n730, Z => n685);
   U1181 : CLKBUF_X1 port map( A => n730, Z => n686);
   U1182 : CLKBUF_X1 port map( A => n730, Z => n687);
   U1183 : CLKBUF_X1 port map( A => n729, Z => n688);
   U1184 : CLKBUF_X1 port map( A => n729, Z => n689);
   U1185 : CLKBUF_X1 port map( A => n729, Z => n690);
   U1186 : CLKBUF_X1 port map( A => n729, Z => n691);
   U1187 : CLKBUF_X1 port map( A => n729, Z => n692);
   U1188 : CLKBUF_X1 port map( A => n728, Z => n693);
   U1189 : CLKBUF_X1 port map( A => n728, Z => n694);
   U1190 : CLKBUF_X1 port map( A => n728, Z => n695);
   U1191 : CLKBUF_X1 port map( A => n728, Z => n696);
   U1192 : CLKBUF_X1 port map( A => n728, Z => n697);
   U1193 : CLKBUF_X1 port map( A => n727, Z => n698);
   U1194 : CLKBUF_X1 port map( A => n727, Z => n699);
   U1195 : CLKBUF_X1 port map( A => n727, Z => n700);
   U1196 : CLKBUF_X1 port map( A => n727, Z => n701);
   U1197 : CLKBUF_X1 port map( A => n727, Z => n702);
   U1198 : CLKBUF_X1 port map( A => n726, Z => n703);
   U1199 : CLKBUF_X1 port map( A => n726, Z => n704);
   U1200 : CLKBUF_X1 port map( A => n726, Z => n705);
   U1201 : CLKBUF_X1 port map( A => n726, Z => n706);
   U1202 : CLKBUF_X1 port map( A => n726, Z => n707);
   U1203 : CLKBUF_X1 port map( A => n725, Z => n708);
   U1204 : CLKBUF_X1 port map( A => n725, Z => n709);
   U1205 : CLKBUF_X1 port map( A => n725, Z => n710);
   U1206 : CLKBUF_X1 port map( A => n725, Z => n711);
   U1207 : CLKBUF_X1 port map( A => n725, Z => n712);
   U1208 : CLKBUF_X1 port map( A => n724, Z => n713);
   U1209 : CLKBUF_X1 port map( A => n724, Z => n714);
   U1210 : CLKBUF_X1 port map( A => n724, Z => n715);
   U1211 : CLKBUF_X1 port map( A => n724, Z => n716);
   U1212 : CLKBUF_X1 port map( A => n724, Z => n717);
   U1213 : CLKBUF_X1 port map( A => n723, Z => n718);
   U1214 : CLKBUF_X1 port map( A => n723, Z => n719);
   U1215 : CLKBUF_X1 port map( A => n723, Z => n720);
   U1216 : CLKBUF_X1 port map( A => n723, Z => n721);
   U1217 : CLKBUF_X1 port map( A => n723, Z => n722);
   U1218 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n732);
   U1219 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n733);
   U1220 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n734);
   U1221 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n735);
   U1222 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n736);
   U1223 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n737);
   U1224 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n738);
   U1225 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n739);
   U1226 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n740);
   U1227 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n741);
   U1228 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n742);
   U1229 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n743);
   U1230 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n744);
   U1231 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n745);
   U1232 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n746);
   U1233 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n747);
   U1234 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n748);
   U1235 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n749);
   U1236 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n750);
   U1237 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n751);
   U1238 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n752);
   U1239 : CLKBUF_X1 port map( A => r3007_A_0_port, Z => n753);
   U1240 : CLKBUF_X1 port map( A => n813, Z => n754);
   U1241 : CLKBUF_X1 port map( A => n813, Z => n755);
   U1242 : CLKBUF_X1 port map( A => n813, Z => n756);
   U1243 : CLKBUF_X1 port map( A => n812, Z => n757);
   U1244 : CLKBUF_X1 port map( A => n812, Z => n758);
   U1245 : CLKBUF_X1 port map( A => n812, Z => n759);
   U1246 : CLKBUF_X1 port map( A => n812, Z => n760);
   U1247 : CLKBUF_X1 port map( A => n812, Z => n761);
   U1248 : CLKBUF_X1 port map( A => n812, Z => n762);
   U1249 : CLKBUF_X1 port map( A => n811, Z => n763);
   U1250 : CLKBUF_X1 port map( A => n811, Z => n764);
   U1251 : CLKBUF_X1 port map( A => n811, Z => n765);
   U1252 : CLKBUF_X1 port map( A => n811, Z => n766);
   U1253 : CLKBUF_X1 port map( A => n811, Z => n767);
   U1254 : CLKBUF_X1 port map( A => n811, Z => n768);
   U1255 : CLKBUF_X1 port map( A => n810, Z => n769);
   U1256 : CLKBUF_X1 port map( A => n810, Z => n770);
   U1257 : CLKBUF_X1 port map( A => n810, Z => n771);
   U1258 : CLKBUF_X1 port map( A => n810, Z => n772);
   U1259 : CLKBUF_X1 port map( A => n810, Z => n773);
   U1260 : CLKBUF_X1 port map( A => n810, Z => n774);
   U1261 : CLKBUF_X1 port map( A => n809, Z => n775);
   U1262 : CLKBUF_X1 port map( A => n809, Z => n776);
   U1263 : CLKBUF_X1 port map( A => n809, Z => n777);
   U1264 : CLKBUF_X1 port map( A => n809, Z => n778);
   U1265 : CLKBUF_X1 port map( A => n809, Z => n779);
   U1266 : CLKBUF_X1 port map( A => n809, Z => n780);
   U1267 : CLKBUF_X1 port map( A => n808, Z => n781);
   U1268 : CLKBUF_X1 port map( A => n808, Z => n782);
   U1269 : CLKBUF_X1 port map( A => n808, Z => n783);
   U1270 : CLKBUF_X1 port map( A => n808, Z => n784);
   U1271 : CLKBUF_X1 port map( A => n808, Z => n785);
   U1272 : CLKBUF_X1 port map( A => n808, Z => n786);
   U1273 : CLKBUF_X1 port map( A => n807, Z => n787);
   U1274 : CLKBUF_X1 port map( A => n807, Z => n788);
   U1275 : CLKBUF_X1 port map( A => n807, Z => n789);
   U1276 : CLKBUF_X1 port map( A => n807, Z => n790);
   U1277 : CLKBUF_X1 port map( A => n807, Z => n791);
   U1278 : CLKBUF_X1 port map( A => n807, Z => n792);
   U1279 : CLKBUF_X1 port map( A => n806, Z => n793);
   U1280 : CLKBUF_X1 port map( A => n806, Z => n794);
   U1281 : CLKBUF_X1 port map( A => n806, Z => n795);
   U1282 : CLKBUF_X1 port map( A => n806, Z => n796);
   U1283 : CLKBUF_X1 port map( A => n806, Z => n797);
   U1284 : CLKBUF_X1 port map( A => n806, Z => n798);
   U1285 : CLKBUF_X1 port map( A => n805, Z => n799);
   U1286 : CLKBUF_X1 port map( A => n805, Z => n800);
   U1287 : CLKBUF_X1 port map( A => n805, Z => n801);
   U1288 : CLKBUF_X1 port map( A => n805, Z => n802);
   U1289 : CLKBUF_X1 port map( A => n805, Z => n803);
   U1290 : CLKBUF_X1 port map( A => n805, Z => n804);
   U1291 : CLKBUF_X1 port map( A => SWP_1_port, Z => n814);
   U1292 : CLKBUF_X1 port map( A => SWP_1_port, Z => n815);
   U1293 : CLKBUF_X1 port map( A => SWP_1_port, Z => n816);
   U1294 : CLKBUF_X1 port map( A => SWP_1_port, Z => n817);
   U1295 : CLKBUF_X1 port map( A => SWP_1_port, Z => n818);
   U1296 : CLKBUF_X1 port map( A => SWP_1_port, Z => n819);
   U1297 : CLKBUF_X1 port map( A => SWP_1_port, Z => n820);
   U1298 : CLKBUF_X1 port map( A => SWP_1_port, Z => n821);
   U1299 : CLKBUF_X1 port map( A => SWP_1_port, Z => n822);
   U1300 : CLKBUF_X1 port map( A => SWP_1_port, Z => n823);
   U1301 : CLKBUF_X1 port map( A => SWP_1_port, Z => n824);
   U1302 : CLKBUF_X1 port map( A => SWP_1_port, Z => n825);
   U1303 : CLKBUF_X1 port map( A => SWP_1_port, Z => n826);
   U1304 : CLKBUF_X1 port map( A => SWP_1_port, Z => n827);
   U1305 : CLKBUF_X1 port map( A => SWP_1_port, Z => n828);
   U1306 : CLKBUF_X1 port map( A => SWP_1_port, Z => n829);
   U1307 : CLKBUF_X1 port map( A => SWP_1_port, Z => n830);
   U1308 : CLKBUF_X1 port map( A => SWP_1_port, Z => n831);
   U1309 : CLKBUF_X1 port map( A => SWP_1_port, Z => n832);
   U1310 : CLKBUF_X1 port map( A => SWP_1_port, Z => n833);
   U1311 : CLKBUF_X1 port map( A => SWP_1_port, Z => n834);
   U1312 : CLKBUF_X1 port map( A => SWP_1_port, Z => n835);
   U1313 : CLKBUF_X1 port map( A => SWP_1_port, Z => n836);
   U1314 : CLKBUF_X1 port map( A => SWP_1_port, Z => n837);
   U1315 : CLKBUF_X1 port map( A => SWP_1_port, Z => n838);
   U1316 : CLKBUF_X1 port map( A => SWP_1_port, Z => n839);
   U1317 : CLKBUF_X1 port map( A => SWP_1_port, Z => n840);
   U1318 : CLKBUF_X1 port map( A => n1003, Z => n850);
   U1319 : CLKBUF_X1 port map( A => n1003, Z => n851);
   U1320 : CLKBUF_X1 port map( A => n1003, Z => n852);
   U1321 : CLKBUF_X1 port map( A => n1003, Z => n853);
   U1322 : CLKBUF_X1 port map( A => n1003, Z => n854);
   U1323 : CLKBUF_X1 port map( A => n1003, Z => n855);
   U1324 : CLKBUF_X1 port map( A => n1002, Z => n856);
   U1325 : CLKBUF_X1 port map( A => n1002, Z => n857);
   U1326 : CLKBUF_X1 port map( A => n1002, Z => n858);
   U1327 : CLKBUF_X1 port map( A => n1002, Z => n859);
   U1328 : CLKBUF_X1 port map( A => n1002, Z => n860);
   U1329 : CLKBUF_X1 port map( A => n1002, Z => n861);
   U1330 : CLKBUF_X1 port map( A => n1001, Z => n862);
   U1331 : CLKBUF_X1 port map( A => n1001, Z => n863);
   U1332 : CLKBUF_X1 port map( A => n1001, Z => n864);
   U1333 : CLKBUF_X1 port map( A => n1001, Z => n865);
   U1334 : CLKBUF_X1 port map( A => n1001, Z => n866);
   U1335 : CLKBUF_X1 port map( A => n1001, Z => n867);
   U1336 : CLKBUF_X1 port map( A => n1000, Z => n868);
   U1337 : CLKBUF_X1 port map( A => n1000, Z => n869);
   U1338 : CLKBUF_X1 port map( A => n1000, Z => n870);
   U1339 : CLKBUF_X1 port map( A => n1000, Z => n871);
   U1340 : CLKBUF_X1 port map( A => n1000, Z => n872);
   U1341 : CLKBUF_X1 port map( A => n1000, Z => n873);
   U1342 : CLKBUF_X1 port map( A => n999, Z => n874);
   U1343 : CLKBUF_X1 port map( A => n999, Z => n875);
   U1344 : CLKBUF_X1 port map( A => n999, Z => n876);
   U1345 : CLKBUF_X1 port map( A => n999, Z => n877);
   U1346 : CLKBUF_X1 port map( A => n999, Z => n878);
   U1347 : CLKBUF_X1 port map( A => n999, Z => n879);
   U1348 : CLKBUF_X1 port map( A => n998, Z => n880);
   U1349 : CLKBUF_X1 port map( A => n998, Z => n881);
   U1350 : CLKBUF_X1 port map( A => n998, Z => n882);
   U1351 : CLKBUF_X1 port map( A => n998, Z => n883);
   U1352 : CLKBUF_X1 port map( A => n998, Z => n884);
   U1353 : CLKBUF_X1 port map( A => n998, Z => n885);
   U1354 : CLKBUF_X1 port map( A => n997, Z => n886);
   U1355 : CLKBUF_X1 port map( A => n997, Z => n887);
   U1356 : CLKBUF_X1 port map( A => n997, Z => n888);
   U1357 : CLKBUF_X1 port map( A => n997, Z => n889);
   U1358 : CLKBUF_X1 port map( A => n997, Z => n890);
   U1359 : CLKBUF_X1 port map( A => n997, Z => n891);
   U1360 : CLKBUF_X1 port map( A => n996, Z => n892);
   U1361 : CLKBUF_X1 port map( A => n996, Z => n893);
   U1362 : CLKBUF_X1 port map( A => n996, Z => n894);
   U1363 : CLKBUF_X1 port map( A => n996, Z => n895);
   U1364 : CLKBUF_X1 port map( A => n996, Z => n896);
   U1365 : CLKBUF_X1 port map( A => n996, Z => n897);
   U1366 : CLKBUF_X1 port map( A => n995, Z => n898);
   U1367 : CLKBUF_X1 port map( A => n995, Z => n899);
   U1368 : CLKBUF_X1 port map( A => n995, Z => n900);
   U1369 : CLKBUF_X1 port map( A => n995, Z => n901);
   U1370 : CLKBUF_X1 port map( A => n995, Z => n902);
   U1371 : CLKBUF_X1 port map( A => n995, Z => n903);
   U1372 : CLKBUF_X1 port map( A => n994, Z => n904);
   U1373 : CLKBUF_X1 port map( A => n994, Z => n905);
   U1374 : CLKBUF_X1 port map( A => n994, Z => n906);
   U1375 : CLKBUF_X1 port map( A => n994, Z => n907);
   U1376 : CLKBUF_X1 port map( A => n994, Z => n908);
   U1377 : CLKBUF_X1 port map( A => n994, Z => n909);
   U1378 : CLKBUF_X1 port map( A => n993, Z => n910);
   U1379 : CLKBUF_X1 port map( A => n993, Z => n911);
   U1380 : CLKBUF_X1 port map( A => n993, Z => n912);
   U1381 : CLKBUF_X1 port map( A => n993, Z => n913);
   U1382 : CLKBUF_X1 port map( A => n993, Z => n914);
   U1383 : CLKBUF_X1 port map( A => n993, Z => n915);
   U1384 : CLKBUF_X1 port map( A => n992, Z => n916);
   U1385 : CLKBUF_X1 port map( A => n992, Z => n917);
   U1386 : CLKBUF_X1 port map( A => n992, Z => n918);
   U1387 : CLKBUF_X1 port map( A => n992, Z => n919);
   U1388 : CLKBUF_X1 port map( A => n992, Z => n920);
   U1389 : CLKBUF_X1 port map( A => n992, Z => n921);
   U1390 : CLKBUF_X1 port map( A => n991, Z => n922);
   U1391 : CLKBUF_X1 port map( A => n991, Z => n923);
   U1392 : CLKBUF_X1 port map( A => n991, Z => n924);
   U1393 : CLKBUF_X1 port map( A => n991, Z => n925);
   U1394 : CLKBUF_X1 port map( A => n991, Z => n926);
   U1395 : CLKBUF_X1 port map( A => n991, Z => n927);
   U1396 : CLKBUF_X1 port map( A => n990, Z => n928);
   U1397 : CLKBUF_X1 port map( A => n990, Z => n929);
   U1398 : CLKBUF_X1 port map( A => n990, Z => n930);
   U1399 : CLKBUF_X1 port map( A => n990, Z => n931);
   U1400 : CLKBUF_X1 port map( A => n990, Z => n932);
   U1401 : CLKBUF_X1 port map( A => n990, Z => n933);
   U1402 : CLKBUF_X1 port map( A => n989, Z => n934);
   U1403 : CLKBUF_X1 port map( A => n989, Z => n935);
   U1404 : CLKBUF_X1 port map( A => n989, Z => n936);
   U1405 : CLKBUF_X1 port map( A => n989, Z => n937);
   U1406 : CLKBUF_X1 port map( A => n989, Z => n938);
   U1407 : CLKBUF_X1 port map( A => n989, Z => n939);
   U1408 : CLKBUF_X1 port map( A => n988, Z => n940);
   U1409 : CLKBUF_X1 port map( A => n988, Z => n941);
   U1410 : CLKBUF_X1 port map( A => n988, Z => n942);
   U1411 : CLKBUF_X1 port map( A => n988, Z => n943);
   U1412 : CLKBUF_X1 port map( A => n988, Z => n944);
   U1413 : CLKBUF_X1 port map( A => n988, Z => n945);
   U1414 : CLKBUF_X1 port map( A => n987, Z => n946);
   U1415 : CLKBUF_X1 port map( A => n987, Z => n947);
   U1416 : CLKBUF_X1 port map( A => n987, Z => n948);
   U1417 : CLKBUF_X1 port map( A => n987, Z => n949);
   U1418 : CLKBUF_X1 port map( A => n987, Z => n950);
   U1419 : CLKBUF_X1 port map( A => n987, Z => n951);
   U1420 : CLKBUF_X1 port map( A => n986, Z => n952);
   U1421 : CLKBUF_X1 port map( A => n986, Z => n953);
   U1422 : CLKBUF_X1 port map( A => n986, Z => n954);
   U1423 : CLKBUF_X1 port map( A => n986, Z => n955);
   U1424 : CLKBUF_X1 port map( A => n986, Z => n956);
   U1425 : CLKBUF_X1 port map( A => n986, Z => n957);
   U1426 : CLKBUF_X1 port map( A => n985, Z => n958);
   U1427 : CLKBUF_X1 port map( A => n985, Z => n959);
   U1428 : CLKBUF_X1 port map( A => n985, Z => n960);
   U1429 : CLKBUF_X1 port map( A => n985, Z => n961);
   U1430 : CLKBUF_X1 port map( A => n985, Z => n962);
   U1431 : CLKBUF_X1 port map( A => n985, Z => n963);
   U1432 : CLKBUF_X1 port map( A => n984, Z => n964);
   U1433 : CLKBUF_X1 port map( A => n984, Z => n965);
   U1434 : CLKBUF_X1 port map( A => n984, Z => n966);
   U1435 : CLKBUF_X1 port map( A => n984, Z => n967);
   U1436 : CLKBUF_X1 port map( A => n984, Z => n968);
   U1437 : CLKBUF_X1 port map( A => n984, Z => n969);
   U1438 : CLKBUF_X1 port map( A => n983, Z => n970);
   U1439 : CLKBUF_X1 port map( A => n983, Z => n971);
   U1440 : CLKBUF_X1 port map( A => n983, Z => n972);
   U1441 : CLKBUF_X1 port map( A => n983, Z => n973);
   U1442 : CLKBUF_X1 port map( A => n983, Z => n974);
   U1443 : CLKBUF_X1 port map( A => n983, Z => n975);
   U1444 : CLKBUF_X1 port map( A => n982, Z => n976);
   U1445 : CLKBUF_X1 port map( A => n982, Z => n977);
   U1446 : CLKBUF_X1 port map( A => n982, Z => n978);
   U1447 : CLKBUF_X1 port map( A => n982, Z => n979);
   U1448 : CLKBUF_X1 port map( A => n982, Z => n980);
   U1449 : CLKBUF_X1 port map( A => n982, Z => n981);
   U1450 : MUX2_X1 port map( A => REGISTERS_5_0_port, B => REGISTERS_6_0_port, 
                           S => n792, Z => n1007);
   U1451 : MUX2_X1 port map( A => REGISTERS_3_0_port, B => REGISTERS_4_0_port, 
                           S => n791, Z => n1008);
   U1452 : MUX2_X1 port map( A => n1008, B => n1007, S => n827, Z => n1009);
   U1453 : MUX2_X1 port map( A => REGISTERS_37_0_port, B => REGISTERS_38_0_port
                           , S => n791, Z => n1010);
   U1454 : MUX2_X1 port map( A => REGISTERS_35_0_port, B => REGISTERS_36_0_port
                           , S => n791, Z => n1011);
   U1455 : MUX2_X1 port map( A => n1011, B => n1010, S => n827, Z => n1012);
   U1456 : MUX2_X1 port map( A => REGISTERS_21_0_port, B => REGISTERS_22_0_port
                           , S => n791, Z => n1013);
   U1457 : MUX2_X1 port map( A => REGISTERS_19_0_port, B => REGISTERS_20_0_port
                           , S => n791, Z => n1014);
   U1458 : MUX2_X1 port map( A => n1014, B => n1013, S => n827, Z => n1015);
   U1459 : MUX2_X1 port map( A => n1015, B => n1012, S => n841, Z => n1016);
   U1460 : MUX2_X1 port map( A => n1016, B => n1009, S => n846, Z => n1017);
   U1461 : MUX2_X1 port map( A => REGISTERS_29_0_port, B => REGISTERS_30_0_port
                           , S => n791, Z => n1018);
   U1462 : MUX2_X1 port map( A => REGISTERS_27_0_port, B => REGISTERS_28_0_port
                           , S => n791, Z => n1019);
   U1463 : MUX2_X1 port map( A => n1019, B => n1018, S => n827, Z => n1020);
   U1464 : MUX2_X1 port map( A => REGISTERS_13_0_port, B => REGISTERS_14_0_port
                           , S => n791, Z => n1021);
   U1465 : MUX2_X1 port map( A => REGISTERS_11_0_port, B => REGISTERS_12_0_port
                           , S => n791, Z => n1022);
   U1466 : MUX2_X1 port map( A => n1022, B => n1021, S => n827, Z => n1023);
   U1467 : MUX2_X1 port map( A => n1023, B => n1020, S => n845, Z => n1024);
   U1468 : MUX2_X1 port map( A => n1024, B => n1017, S => n302, Z => n1025);
   U1469 : MUX2_X1 port map( A => REGISTERS_1_0_port, B => REGISTERS_2_0_port, 
                           S => n791, Z => n1026);
   U1470 : MUX2_X1 port map( A => REGISTERS_0_0_port, B => n1026, S => n827, Z 
                           => n1027);
   U1471 : MUX2_X1 port map( A => REGISTERS_33_0_port, B => REGISTERS_34_0_port
                           , S => n791, Z => n1028);
   U1472 : MUX2_X1 port map( A => REGISTERS_31_0_port, B => REGISTERS_32_0_port
                           , S => n791, Z => n1029);
   U1473 : MUX2_X1 port map( A => n1029, B => n1028, S => n828, Z => n1030);
   U1474 : MUX2_X1 port map( A => REGISTERS_17_0_port, B => REGISTERS_18_0_port
                           , S => n790, Z => n1031);
   U1475 : MUX2_X1 port map( A => REGISTERS_15_0_port, B => REGISTERS_16_0_port
                           , S => n790, Z => n1032);
   U1476 : MUX2_X1 port map( A => n1032, B => n1031, S => n828, Z => n1033);
   U1477 : MUX2_X1 port map( A => n1033, B => n1030, S => n845, Z => n1034);
   U1478 : MUX2_X1 port map( A => n1034, B => n1027, S => n849, Z => n1035);
   U1479 : MUX2_X1 port map( A => REGISTERS_25_0_port, B => REGISTERS_26_0_port
                           , S => n790, Z => n1036);
   U1480 : MUX2_X1 port map( A => REGISTERS_23_0_port, B => REGISTERS_24_0_port
                           , S => n790, Z => n1037);
   U1481 : MUX2_X1 port map( A => n1037, B => n1036, S => n828, Z => n1038);
   U1482 : MUX2_X1 port map( A => REGISTERS_9_0_port, B => REGISTERS_10_0_port,
                           S => n790, Z => n1039);
   U1483 : MUX2_X1 port map( A => REGISTERS_7_0_port, B => REGISTERS_8_0_port, 
                           S => n790, Z => n1040);
   U1484 : MUX2_X1 port map( A => n1040, B => n1039, S => n828, Z => n1041);
   U1485 : MUX2_X1 port map( A => n1041, B => n1038, S => n845, Z => n1042);
   U1486 : MUX2_X1 port map( A => n1042, B => REGISTERS_39_0_port, S => n849, Z
                           => n1043);
   U1487 : MUX2_X1 port map( A => n1043, B => n1035, S => n302, Z => n1044);
   U1488 : MUX2_X1 port map( A => n1044, B => n1025, S => n301, Z => N12205);
   U1489 : MUX2_X1 port map( A => REGISTERS_5_1_port, B => REGISTERS_6_1_port, 
                           S => n790, Z => n1045);
   U1490 : MUX2_X1 port map( A => REGISTERS_3_1_port, B => REGISTERS_4_1_port, 
                           S => n790, Z => n1046);
   U1491 : MUX2_X1 port map( A => n1046, B => n1045, S => n828, Z => n1047);
   U1492 : MUX2_X1 port map( A => REGISTERS_37_1_port, B => REGISTERS_38_1_port
                           , S => n790, Z => n1048);
   U1493 : MUX2_X1 port map( A => REGISTERS_35_1_port, B => REGISTERS_36_1_port
                           , S => n790, Z => n1049);
   U1494 : MUX2_X1 port map( A => n1049, B => n1048, S => n828, Z => n1050);
   U1495 : MUX2_X1 port map( A => REGISTERS_21_1_port, B => REGISTERS_22_1_port
                           , S => n790, Z => n1051);
   U1496 : MUX2_X1 port map( A => REGISTERS_19_1_port, B => REGISTERS_20_1_port
                           , S => n790, Z => n1052);
   U1497 : MUX2_X1 port map( A => n1052, B => n1051, S => n828, Z => n1053);
   U1498 : MUX2_X1 port map( A => n1053, B => n1050, S => n845, Z => n1054);
   U1499 : MUX2_X1 port map( A => n1054, B => n1047, S => n849, Z => n1055);
   U1500 : MUX2_X1 port map( A => REGISTERS_29_1_port, B => REGISTERS_30_1_port
                           , S => n789, Z => n1056);
   U1501 : MUX2_X1 port map( A => REGISTERS_27_1_port, B => REGISTERS_28_1_port
                           , S => n789, Z => n1057);
   U1502 : MUX2_X1 port map( A => n1057, B => n1056, S => n828, Z => n1058);
   U1503 : MUX2_X1 port map( A => REGISTERS_13_1_port, B => REGISTERS_14_1_port
                           , S => n789, Z => n1059);
   U1504 : MUX2_X1 port map( A => REGISTERS_11_1_port, B => REGISTERS_12_1_port
                           , S => n789, Z => n1060);
   U1505 : MUX2_X1 port map( A => n1060, B => n1059, S => n828, Z => n1061);
   U1506 : MUX2_X1 port map( A => n1061, B => n1058, S => n845, Z => n1062);
   U1507 : MUX2_X1 port map( A => n1062, B => n1055, S => n302, Z => n1063);
   U1508 : MUX2_X1 port map( A => REGISTERS_1_1_port, B => REGISTERS_2_1_port, 
                           S => n789, Z => n1064);
   U1509 : MUX2_X1 port map( A => REGISTERS_0_1_port, B => n1064, S => n828, Z 
                           => n1065);
   U1510 : MUX2_X1 port map( A => REGISTERS_33_1_port, B => REGISTERS_34_1_port
                           , S => n789, Z => n1066);
   U1511 : MUX2_X1 port map( A => REGISTERS_31_1_port, B => REGISTERS_32_1_port
                           , S => n789, Z => n1067);
   U1512 : MUX2_X1 port map( A => n1067, B => n1066, S => n828, Z => n1068);
   U1513 : MUX2_X1 port map( A => REGISTERS_17_1_port, B => REGISTERS_18_1_port
                           , S => n789, Z => n1069);
   U1514 : MUX2_X1 port map( A => REGISTERS_15_1_port, B => REGISTERS_16_1_port
                           , S => n789, Z => n1070);
   U1515 : MUX2_X1 port map( A => n1070, B => n1069, S => n828, Z => n1071);
   U1516 : MUX2_X1 port map( A => n1071, B => n1068, S => n845, Z => n1072);
   U1517 : MUX2_X1 port map( A => n1072, B => n1065, S => n849, Z => n1073);
   U1518 : MUX2_X1 port map( A => REGISTERS_25_1_port, B => REGISTERS_26_1_port
                           , S => n789, Z => n1074);
   U1519 : MUX2_X1 port map( A => REGISTERS_23_1_port, B => REGISTERS_24_1_port
                           , S => n789, Z => n1075);
   U1520 : MUX2_X1 port map( A => n1075, B => n1074, S => n829, Z => n1076);
   U1521 : MUX2_X1 port map( A => REGISTERS_9_1_port, B => REGISTERS_10_1_port,
                           S => n789, Z => n1077);
   U1522 : MUX2_X1 port map( A => REGISTERS_7_1_port, B => REGISTERS_8_1_port, 
                           S => n788, Z => n1078);
   U1523 : MUX2_X1 port map( A => n1078, B => n1077, S => n829, Z => n1079);
   U1524 : MUX2_X1 port map( A => n1079, B => n1076, S => n845, Z => n1080);
   U1525 : MUX2_X1 port map( A => n1080, B => REGISTERS_39_1_port, S => n849, Z
                           => n1081);
   U1526 : MUX2_X1 port map( A => n1081, B => n1073, S => n302, Z => n1082);
   U1527 : MUX2_X1 port map( A => n1082, B => n1063, S => n301, Z => N12206);
   U1528 : MUX2_X1 port map( A => REGISTERS_5_2_port, B => REGISTERS_6_2_port, 
                           S => n788, Z => n1083);
   U1529 : MUX2_X1 port map( A => REGISTERS_3_2_port, B => REGISTERS_4_2_port, 
                           S => n788, Z => n1084);
   U1530 : MUX2_X1 port map( A => n1084, B => n1083, S => n829, Z => n1085);
   U1531 : MUX2_X1 port map( A => REGISTERS_37_2_port, B => REGISTERS_38_2_port
                           , S => n788, Z => n1086);
   U1532 : MUX2_X1 port map( A => REGISTERS_35_2_port, B => REGISTERS_36_2_port
                           , S => n788, Z => n1087);
   U1533 : MUX2_X1 port map( A => n1087, B => n1086, S => n829, Z => n1088);
   U1534 : MUX2_X1 port map( A => REGISTERS_21_2_port, B => REGISTERS_22_2_port
                           , S => n788, Z => n1089);
   U1535 : MUX2_X1 port map( A => REGISTERS_19_2_port, B => REGISTERS_20_2_port
                           , S => n788, Z => n1090);
   U1536 : MUX2_X1 port map( A => n1090, B => n1089, S => n829, Z => n1091);
   U1537 : MUX2_X1 port map( A => n1091, B => n1088, S => n845, Z => n1092);
   U1538 : MUX2_X1 port map( A => n1092, B => n1085, S => n849, Z => n1093);
   U1539 : MUX2_X1 port map( A => REGISTERS_29_2_port, B => REGISTERS_30_2_port
                           , S => n788, Z => n1094);
   U1540 : MUX2_X1 port map( A => REGISTERS_27_2_port, B => REGISTERS_28_2_port
                           , S => n788, Z => n1095);
   U1541 : MUX2_X1 port map( A => n1095, B => n1094, S => n829, Z => n1096);
   U1542 : MUX2_X1 port map( A => REGISTERS_13_2_port, B => REGISTERS_14_2_port
                           , S => n788, Z => n1097);
   U1543 : MUX2_X1 port map( A => REGISTERS_11_2_port, B => REGISTERS_12_2_port
                           , S => n788, Z => n1098);
   U1544 : MUX2_X1 port map( A => n1098, B => n1097, S => n829, Z => n1099);
   U1545 : MUX2_X1 port map( A => n1099, B => n1096, S => n845, Z => n1100);
   U1546 : MUX2_X1 port map( A => n1100, B => n1093, S => n302, Z => n1101);
   U1547 : MUX2_X1 port map( A => REGISTERS_1_2_port, B => REGISTERS_2_2_port, 
                           S => n788, Z => n1102);
   U1548 : MUX2_X1 port map( A => REGISTERS_0_2_port, B => n1102, S => n829, Z 
                           => n1103);
   U1549 : MUX2_X1 port map( A => REGISTERS_33_2_port, B => REGISTERS_34_2_port
                           , S => n787, Z => n1104);
   U1550 : MUX2_X1 port map( A => REGISTERS_31_2_port, B => REGISTERS_32_2_port
                           , S => n787, Z => n1105);
   U1551 : MUX2_X1 port map( A => n1105, B => n1104, S => n829, Z => n1106);
   U1552 : MUX2_X1 port map( A => REGISTERS_17_2_port, B => REGISTERS_18_2_port
                           , S => n787, Z => n1107);
   U1553 : MUX2_X1 port map( A => REGISTERS_15_2_port, B => REGISTERS_16_2_port
                           , S => n787, Z => n1108);
   U1554 : MUX2_X1 port map( A => n1108, B => n1107, S => n829, Z => n1109);
   U1555 : MUX2_X1 port map( A => n1109, B => n1106, S => n845, Z => n1110);
   U1556 : MUX2_X1 port map( A => n1110, B => n1103, S => n849, Z => n1111);
   U1557 : MUX2_X1 port map( A => REGISTERS_25_2_port, B => REGISTERS_26_2_port
                           , S => n787, Z => n1112);
   U1558 : MUX2_X1 port map( A => REGISTERS_23_2_port, B => REGISTERS_24_2_port
                           , S => n787, Z => n1113);
   U1559 : MUX2_X1 port map( A => n1113, B => n1112, S => n829, Z => n1114);
   U1560 : MUX2_X1 port map( A => REGISTERS_9_2_port, B => REGISTERS_10_2_port,
                           S => n787, Z => n1115);
   U1561 : MUX2_X1 port map( A => REGISTERS_7_2_port, B => REGISTERS_8_2_port, 
                           S => n787, Z => n1116);
   U1562 : MUX2_X1 port map( A => n1116, B => n1115, S => n829, Z => n1117);
   U1563 : MUX2_X1 port map( A => n1117, B => n1114, S => n845, Z => n1118);
   U1564 : MUX2_X1 port map( A => n1118, B => REGISTERS_39_2_port, S => n849, Z
                           => n1119);
   U1565 : MUX2_X1 port map( A => n1119, B => n1111, S => n302, Z => n1120);
   U1566 : MUX2_X1 port map( A => n1120, B => n1101, S => n301, Z => N12207);
   U1567 : MUX2_X1 port map( A => REGISTERS_5_3_port, B => REGISTERS_6_3_port, 
                           S => n787, Z => n1121);
   U1568 : MUX2_X1 port map( A => REGISTERS_3_3_port, B => REGISTERS_4_3_port, 
                           S => n787, Z => n1122);
   U1569 : MUX2_X1 port map( A => n1122, B => n1121, S => n830, Z => n1123);
   U1570 : MUX2_X1 port map( A => REGISTERS_37_3_port, B => REGISTERS_38_3_port
                           , S => n787, Z => n1124);
   U1571 : MUX2_X1 port map( A => REGISTERS_35_3_port, B => REGISTERS_36_3_port
                           , S => n787, Z => n1125);
   U1572 : MUX2_X1 port map( A => n1125, B => n1124, S => n830, Z => n1126);
   U1573 : MUX2_X1 port map( A => REGISTERS_21_3_port, B => REGISTERS_22_3_port
                           , S => n786, Z => n1127);
   U1574 : MUX2_X1 port map( A => REGISTERS_19_3_port, B => REGISTERS_20_3_port
                           , S => n786, Z => n1128);
   U1575 : MUX2_X1 port map( A => n1128, B => n1127, S => n830, Z => n1129);
   U1576 : MUX2_X1 port map( A => n1129, B => n1126, S => n845, Z => n1130);
   U1577 : MUX2_X1 port map( A => n1130, B => n1123, S => n849, Z => n1131);
   U1578 : MUX2_X1 port map( A => REGISTERS_29_3_port, B => REGISTERS_30_3_port
                           , S => n786, Z => n1132);
   U1579 : MUX2_X1 port map( A => REGISTERS_27_3_port, B => REGISTERS_28_3_port
                           , S => n786, Z => n1133);
   U1580 : MUX2_X1 port map( A => n1133, B => n1132, S => n830, Z => n1134);
   U1581 : MUX2_X1 port map( A => REGISTERS_13_3_port, B => REGISTERS_14_3_port
                           , S => n786, Z => n1135);
   U1582 : MUX2_X1 port map( A => REGISTERS_11_3_port, B => REGISTERS_12_3_port
                           , S => n786, Z => n1136);
   U1583 : MUX2_X1 port map( A => n1136, B => n1135, S => n830, Z => n1137);
   U1584 : MUX2_X1 port map( A => n1137, B => n1134, S => n845, Z => n1138);
   U1585 : MUX2_X1 port map( A => n1138, B => n1131, S => n302, Z => n1139);
   U1586 : MUX2_X1 port map( A => REGISTERS_1_3_port, B => REGISTERS_2_3_port, 
                           S => n786, Z => n1140);
   U1587 : MUX2_X1 port map( A => REGISTERS_0_3_port, B => n1140, S => n830, Z 
                           => n1141);
   U1588 : MUX2_X1 port map( A => REGISTERS_33_3_port, B => REGISTERS_34_3_port
                           , S => n786, Z => n1142);
   U1589 : MUX2_X1 port map( A => REGISTERS_31_3_port, B => REGISTERS_32_3_port
                           , S => n786, Z => n1143);
   U1590 : MUX2_X1 port map( A => n1143, B => n1142, S => n830, Z => n1144);
   U1591 : MUX2_X1 port map( A => REGISTERS_17_3_port, B => REGISTERS_18_3_port
                           , S => n786, Z => n1145);
   U1592 : MUX2_X1 port map( A => REGISTERS_15_3_port, B => REGISTERS_16_3_port
                           , S => n786, Z => n1146);
   U1593 : MUX2_X1 port map( A => n1146, B => n1145, S => n830, Z => n1147);
   U1594 : MUX2_X1 port map( A => n1147, B => n1144, S => n845, Z => n1148);
   U1595 : MUX2_X1 port map( A => n1148, B => n1141, S => n849, Z => n1149);
   U1596 : MUX2_X1 port map( A => REGISTERS_25_3_port, B => REGISTERS_26_3_port
                           , S => n786, Z => n1150);
   U1597 : MUX2_X1 port map( A => REGISTERS_23_3_port, B => REGISTERS_24_3_port
                           , S => n785, Z => n1151);
   U1598 : MUX2_X1 port map( A => n1151, B => n1150, S => n830, Z => n1152);
   U1599 : MUX2_X1 port map( A => REGISTERS_9_3_port, B => REGISTERS_10_3_port,
                           S => n785, Z => n1153);
   U1600 : MUX2_X1 port map( A => REGISTERS_7_3_port, B => REGISTERS_8_3_port, 
                           S => n792, Z => n1154);
   U1601 : MUX2_X1 port map( A => n1154, B => n1153, S => n834, Z => n1155);
   U1602 : MUX2_X1 port map( A => n1155, B => n1152, S => n845, Z => n1156);
   U1603 : MUX2_X1 port map( A => n1156, B => REGISTERS_39_3_port, S => n849, Z
                           => n1157);
   U1604 : MUX2_X1 port map( A => n1157, B => n1149, S => n302, Z => n1158);
   U1605 : MUX2_X1 port map( A => n1158, B => n1139, S => n301, Z => N12208);
   U1606 : MUX2_X1 port map( A => REGISTERS_5_4_port, B => REGISTERS_6_4_port, 
                           S => n785, Z => n1159);
   U1607 : MUX2_X1 port map( A => REGISTERS_3_4_port, B => REGISTERS_4_4_port, 
                           S => n785, Z => n1160);
   U1608 : MUX2_X1 port map( A => n1160, B => n1159, S => n830, Z => n1161);
   U1609 : MUX2_X1 port map( A => REGISTERS_37_4_port, B => REGISTERS_38_4_port
                           , S => n785, Z => n1162);
   U1610 : MUX2_X1 port map( A => REGISTERS_35_4_port, B => REGISTERS_36_4_port
                           , S => n785, Z => n1163);
   U1611 : MUX2_X1 port map( A => n1163, B => n1162, S => n830, Z => n1164);
   U1612 : MUX2_X1 port map( A => REGISTERS_21_4_port, B => REGISTERS_22_4_port
                           , S => n785, Z => n1165);
   U1613 : MUX2_X1 port map( A => REGISTERS_19_4_port, B => REGISTERS_20_4_port
                           , S => n785, Z => n1166);
   U1614 : MUX2_X1 port map( A => n1166, B => n1165, S => n830, Z => n1167);
   U1615 : MUX2_X1 port map( A => n1167, B => n1164, S => n845, Z => n1168);
   U1616 : MUX2_X1 port map( A => n1168, B => n1161, S => n849, Z => n1169);
   U1617 : MUX2_X1 port map( A => REGISTERS_29_4_port, B => REGISTERS_30_4_port
                           , S => n785, Z => n1170);
   U1618 : MUX2_X1 port map( A => REGISTERS_27_4_port, B => REGISTERS_28_4_port
                           , S => n785, Z => n1171);
   U1619 : MUX2_X1 port map( A => n1171, B => n1170, S => n831, Z => n1172);
   U1620 : MUX2_X1 port map( A => REGISTERS_13_4_port, B => REGISTERS_14_4_port
                           , S => n785, Z => n1173);
   U1621 : MUX2_X1 port map( A => REGISTERS_11_4_port, B => REGISTERS_12_4_port
                           , S => n784, Z => n1174);
   U1622 : MUX2_X1 port map( A => n1174, B => n1173, S => n831, Z => n1175);
   U1623 : MUX2_X1 port map( A => n1175, B => n1172, S => n844, Z => n1176);
   U1624 : MUX2_X1 port map( A => n1176, B => n1169, S => n302, Z => n1177);
   U1625 : MUX2_X1 port map( A => REGISTERS_1_4_port, B => REGISTERS_2_4_port, 
                           S => n784, Z => n1178);
   U1626 : MUX2_X1 port map( A => REGISTERS_0_4_port, B => n1178, S => n831, Z 
                           => n1179);
   U1627 : MUX2_X1 port map( A => REGISTERS_33_4_port, B => REGISTERS_34_4_port
                           , S => n784, Z => n1180);
   U1628 : MUX2_X1 port map( A => REGISTERS_31_4_port, B => REGISTERS_32_4_port
                           , S => n784, Z => n1181);
   U1629 : MUX2_X1 port map( A => n1181, B => n1180, S => n831, Z => n1182);
   U1630 : MUX2_X1 port map( A => REGISTERS_17_4_port, B => REGISTERS_18_4_port
                           , S => n784, Z => n1183);
   U1631 : MUX2_X1 port map( A => REGISTERS_15_4_port, B => REGISTERS_16_4_port
                           , S => n784, Z => n1184);
   U1632 : MUX2_X1 port map( A => n1184, B => n1183, S => n831, Z => n1185);
   U1633 : MUX2_X1 port map( A => n1185, B => n1182, S => n844, Z => n1186);
   U1634 : MUX2_X1 port map( A => n1186, B => n1179, S => n849, Z => n1187);
   U1635 : MUX2_X1 port map( A => REGISTERS_25_4_port, B => REGISTERS_26_4_port
                           , S => n784, Z => n1188);
   U1636 : MUX2_X1 port map( A => REGISTERS_23_4_port, B => REGISTERS_24_4_port
                           , S => n784, Z => n1189);
   U1637 : MUX2_X1 port map( A => n1189, B => n1188, S => n831, Z => n1190);
   U1638 : MUX2_X1 port map( A => REGISTERS_9_4_port, B => REGISTERS_10_4_port,
                           S => n784, Z => n1191);
   U1639 : MUX2_X1 port map( A => REGISTERS_7_4_port, B => REGISTERS_8_4_port, 
                           S => n784, Z => n1192);
   U1640 : MUX2_X1 port map( A => n1192, B => n1191, S => n831, Z => n1193);
   U1641 : MUX2_X1 port map( A => n1193, B => n1190, S => n844, Z => n1194);
   U1642 : MUX2_X1 port map( A => n1194, B => REGISTERS_39_4_port, S => n849, Z
                           => n1195);
   U1643 : MUX2_X1 port map( A => n1195, B => n1187, S => n302, Z => n1196);
   U1644 : MUX2_X1 port map( A => n1196, B => n1177, S => n301, Z => N12209);
   U1645 : MUX2_X1 port map( A => REGISTERS_5_5_port, B => REGISTERS_6_5_port, 
                           S => n784, Z => n1197);
   U1646 : MUX2_X1 port map( A => REGISTERS_3_5_port, B => REGISTERS_4_5_port, 
                           S => n784, Z => n1198);
   U1647 : MUX2_X1 port map( A => n1198, B => n1197, S => n831, Z => n1199);
   U1648 : MUX2_X1 port map( A => REGISTERS_37_5_port, B => REGISTERS_38_5_port
                           , S => n783, Z => n1200);
   U1649 : MUX2_X1 port map( A => REGISTERS_35_5_port, B => REGISTERS_36_5_port
                           , S => n783, Z => n1201);
   U1650 : MUX2_X1 port map( A => n1201, B => n1200, S => n831, Z => n1202);
   U1651 : MUX2_X1 port map( A => REGISTERS_21_5_port, B => REGISTERS_22_5_port
                           , S => n783, Z => n1203);
   U1652 : MUX2_X1 port map( A => REGISTERS_19_5_port, B => REGISTERS_20_5_port
                           , S => n783, Z => n1204);
   U1653 : MUX2_X1 port map( A => n1204, B => n1203, S => n831, Z => n1205);
   U1654 : MUX2_X1 port map( A => n1205, B => n1202, S => n844, Z => n1206);
   U1655 : MUX2_X1 port map( A => n1206, B => n1199, S => n849, Z => n1207);
   U1656 : MUX2_X1 port map( A => REGISTERS_29_5_port, B => REGISTERS_30_5_port
                           , S => n783, Z => n1208);
   U1657 : MUX2_X1 port map( A => REGISTERS_27_5_port, B => REGISTERS_28_5_port
                           , S => n783, Z => n1209);
   U1658 : MUX2_X1 port map( A => n1209, B => n1208, S => n831, Z => n1210);
   U1659 : MUX2_X1 port map( A => REGISTERS_13_5_port, B => REGISTERS_14_5_port
                           , S => n783, Z => n1211);
   U1660 : MUX2_X1 port map( A => REGISTERS_11_5_port, B => REGISTERS_12_5_port
                           , S => n783, Z => n1212);
   U1661 : MUX2_X1 port map( A => n1212, B => n1211, S => n831, Z => n1213);
   U1662 : MUX2_X1 port map( A => n1213, B => n1210, S => n844, Z => n1214);
   U1663 : MUX2_X1 port map( A => n1214, B => n1207, S => n302, Z => n1215);
   U1664 : MUX2_X1 port map( A => REGISTERS_1_5_port, B => REGISTERS_2_5_port, 
                           S => n783, Z => n1216);
   U1665 : MUX2_X1 port map( A => REGISTERS_0_5_port, B => n1216, S => n832, Z 
                           => n1217);
   U1666 : MUX2_X1 port map( A => REGISTERS_33_5_port, B => REGISTERS_34_5_port
                           , S => n783, Z => n1218);
   U1667 : MUX2_X1 port map( A => REGISTERS_31_5_port, B => REGISTERS_32_5_port
                           , S => n783, Z => n1219);
   U1668 : MUX2_X1 port map( A => n1219, B => n1218, S => n832, Z => n1220);
   U1669 : MUX2_X1 port map( A => REGISTERS_17_5_port, B => REGISTERS_18_5_port
                           , S => n783, Z => n1221);
   U1670 : MUX2_X1 port map( A => REGISTERS_15_5_port, B => REGISTERS_16_5_port
                           , S => n782, Z => n1222);
   U1671 : MUX2_X1 port map( A => n1222, B => n1221, S => n832, Z => n1223);
   U1672 : MUX2_X1 port map( A => n1223, B => n1220, S => n844, Z => n1224);
   U1673 : MUX2_X1 port map( A => n1224, B => n1217, S => n849, Z => n1225);
   U1674 : MUX2_X1 port map( A => REGISTERS_25_5_port, B => REGISTERS_26_5_port
                           , S => n782, Z => n1226);
   U1675 : MUX2_X1 port map( A => REGISTERS_23_5_port, B => REGISTERS_24_5_port
                           , S => n782, Z => n1227);
   U1676 : MUX2_X1 port map( A => n1227, B => n1226, S => n832, Z => n1228);
   U1677 : MUX2_X1 port map( A => REGISTERS_9_5_port, B => REGISTERS_10_5_port,
                           S => n782, Z => n1229);
   U1678 : MUX2_X1 port map( A => REGISTERS_7_5_port, B => REGISTERS_8_5_port, 
                           S => n782, Z => n1230);
   U1679 : MUX2_X1 port map( A => n1230, B => n1229, S => n832, Z => n1231);
   U1680 : MUX2_X1 port map( A => n1231, B => n1228, S => n844, Z => n1232);
   U1681 : MUX2_X1 port map( A => n1232, B => REGISTERS_39_5_port, S => n849, Z
                           => n1233);
   U1682 : MUX2_X1 port map( A => n1233, B => n1225, S => n302, Z => n1234);
   U1683 : MUX2_X1 port map( A => n1234, B => n1215, S => n301, Z => N12210);
   U1684 : MUX2_X1 port map( A => REGISTERS_5_6_port, B => REGISTERS_6_6_port, 
                           S => n782, Z => n1235);
   U1685 : MUX2_X1 port map( A => REGISTERS_3_6_port, B => REGISTERS_4_6_port, 
                           S => n782, Z => n1236);
   U1686 : MUX2_X1 port map( A => n1236, B => n1235, S => n832, Z => n1237);
   U1687 : MUX2_X1 port map( A => REGISTERS_37_6_port, B => REGISTERS_38_6_port
                           , S => n782, Z => n1238);
   U1688 : MUX2_X1 port map( A => REGISTERS_35_6_port, B => REGISTERS_36_6_port
                           , S => n782, Z => n1239);
   U1689 : MUX2_X1 port map( A => n1239, B => n1238, S => n832, Z => n1240);
   U1690 : MUX2_X1 port map( A => REGISTERS_21_6_port, B => REGISTERS_22_6_port
                           , S => n782, Z => n1241);
   U1691 : MUX2_X1 port map( A => REGISTERS_19_6_port, B => REGISTERS_20_6_port
                           , S => n782, Z => n1242);
   U1692 : MUX2_X1 port map( A => n1242, B => n1241, S => n832, Z => n1243);
   U1693 : MUX2_X1 port map( A => n1243, B => n1240, S => n844, Z => n1244);
   U1694 : MUX2_X1 port map( A => n1244, B => n1237, S => n849, Z => n1245);
   U1695 : MUX2_X1 port map( A => REGISTERS_29_6_port, B => REGISTERS_30_6_port
                           , S => n782, Z => n1246);
   U1696 : MUX2_X1 port map( A => REGISTERS_27_6_port, B => REGISTERS_28_6_port
                           , S => n781, Z => n1247);
   U1697 : MUX2_X1 port map( A => n1247, B => n1246, S => n832, Z => n1248);
   U1698 : MUX2_X1 port map( A => REGISTERS_13_6_port, B => REGISTERS_14_6_port
                           , S => n781, Z => n1249);
   U1699 : MUX2_X1 port map( A => REGISTERS_11_6_port, B => REGISTERS_12_6_port
                           , S => n781, Z => n1250);
   U1700 : MUX2_X1 port map( A => n1250, B => n1249, S => n832, Z => n1251);
   U1701 : MUX2_X1 port map( A => n1251, B => n1248, S => n844, Z => n1252);
   U1702 : MUX2_X1 port map( A => n1252, B => n1245, S => n302, Z => n1253);
   U1703 : MUX2_X1 port map( A => REGISTERS_1_6_port, B => REGISTERS_2_6_port, 
                           S => n781, Z => n1254);
   U1704 : MUX2_X1 port map( A => REGISTERS_0_6_port, B => n1254, S => n832, Z 
                           => n1255);
   U1705 : MUX2_X1 port map( A => REGISTERS_33_6_port, B => REGISTERS_34_6_port
                           , S => n781, Z => n1256);
   U1706 : MUX2_X1 port map( A => REGISTERS_31_6_port, B => REGISTERS_32_6_port
                           , S => n781, Z => n1257);
   U1707 : MUX2_X1 port map( A => n1257, B => n1256, S => n832, Z => n1258);
   U1708 : MUX2_X1 port map( A => REGISTERS_17_6_port, B => REGISTERS_18_6_port
                           , S => n781, Z => n1259);
   U1709 : MUX2_X1 port map( A => REGISTERS_15_6_port, B => REGISTERS_16_6_port
                           , S => n781, Z => n1260);
   U1710 : MUX2_X1 port map( A => n1260, B => n1259, S => n833, Z => n1261);
   U1711 : MUX2_X1 port map( A => n1261, B => n1258, S => n844, Z => n1262);
   U1712 : MUX2_X1 port map( A => n1262, B => n1255, S => n849, Z => n1263);
   U1713 : MUX2_X1 port map( A => REGISTERS_25_6_port, B => REGISTERS_26_6_port
                           , S => n781, Z => n1264);
   U1714 : MUX2_X1 port map( A => REGISTERS_23_6_port, B => REGISTERS_24_6_port
                           , S => n781, Z => n1265);
   U1715 : MUX2_X1 port map( A => n1265, B => n1264, S => n833, Z => n1266);
   U1716 : MUX2_X1 port map( A => REGISTERS_9_6_port, B => REGISTERS_10_6_port,
                           S => n781, Z => n1267);
   U1717 : MUX2_X1 port map( A => REGISTERS_7_6_port, B => REGISTERS_8_6_port, 
                           S => n781, Z => n1268);
   U1718 : MUX2_X1 port map( A => n1268, B => n1267, S => n833, Z => n1269);
   U1719 : MUX2_X1 port map( A => n1269, B => n1266, S => n844, Z => n1270);
   U1720 : MUX2_X1 port map( A => n1270, B => REGISTERS_39_6_port, S => n849, Z
                           => n1271);
   U1721 : MUX2_X1 port map( A => n1271, B => n1263, S => n302, Z => n1272);
   U1722 : MUX2_X1 port map( A => n1272, B => n1253, S => n301, Z => N12211);
   U1723 : MUX2_X1 port map( A => REGISTERS_5_7_port, B => REGISTERS_6_7_port, 
                           S => n780, Z => n1273);
   U1724 : MUX2_X1 port map( A => REGISTERS_3_7_port, B => REGISTERS_4_7_port, 
                           S => n780, Z => n1274);
   U1725 : MUX2_X1 port map( A => n1274, B => n1273, S => n833, Z => n1275);
   U1726 : MUX2_X1 port map( A => REGISTERS_37_7_port, B => REGISTERS_38_7_port
                           , S => n780, Z => n1276);
   U1727 : MUX2_X1 port map( A => REGISTERS_35_7_port, B => REGISTERS_36_7_port
                           , S => n780, Z => n1277);
   U1728 : MUX2_X1 port map( A => n1277, B => n1276, S => n833, Z => n1278);
   U1729 : MUX2_X1 port map( A => REGISTERS_21_7_port, B => REGISTERS_22_7_port
                           , S => n780, Z => n1279);
   U1730 : MUX2_X1 port map( A => REGISTERS_19_7_port, B => REGISTERS_20_7_port
                           , S => n780, Z => n1280);
   U1731 : MUX2_X1 port map( A => n1280, B => n1279, S => n833, Z => n1281);
   U1732 : MUX2_X1 port map( A => n1281, B => n1278, S => n844, Z => n1282);
   U1733 : MUX2_X1 port map( A => n1282, B => n1275, S => n849, Z => n1283);
   U1734 : MUX2_X1 port map( A => REGISTERS_29_7_port, B => REGISTERS_30_7_port
                           , S => n780, Z => n1284);
   U1735 : MUX2_X1 port map( A => REGISTERS_27_7_port, B => REGISTERS_28_7_port
                           , S => n780, Z => n1285);
   U1736 : MUX2_X1 port map( A => n1285, B => n1284, S => n833, Z => n1286);
   U1737 : MUX2_X1 port map( A => REGISTERS_13_7_port, B => REGISTERS_14_7_port
                           , S => n780, Z => n1287);
   U1738 : MUX2_X1 port map( A => REGISTERS_11_7_port, B => REGISTERS_12_7_port
                           , S => n780, Z => n1288);
   U1739 : MUX2_X1 port map( A => n1288, B => n1287, S => n833, Z => n1289);
   U1740 : MUX2_X1 port map( A => n1289, B => n1286, S => n844, Z => n1290);
   U1741 : MUX2_X1 port map( A => n1290, B => n1283, S => n302, Z => n1291);
   U1742 : MUX2_X1 port map( A => REGISTERS_1_7_port, B => REGISTERS_2_7_port, 
                           S => n780, Z => n1292);
   U1743 : MUX2_X1 port map( A => REGISTERS_0_7_port, B => n1292, S => n833, Z 
                           => n1293);
   U1744 : MUX2_X1 port map( A => REGISTERS_33_7_port, B => REGISTERS_34_7_port
                           , S => n780, Z => n1294);
   U1745 : MUX2_X1 port map( A => REGISTERS_31_7_port, B => REGISTERS_32_7_port
                           , S => n779, Z => n1295);
   U1746 : MUX2_X1 port map( A => n1295, B => n1294, S => n833, Z => n1296);
   U1747 : MUX2_X1 port map( A => REGISTERS_17_7_port, B => REGISTERS_18_7_port
                           , S => n779, Z => n1297);
   U1748 : MUX2_X1 port map( A => REGISTERS_15_7_port, B => REGISTERS_16_7_port
                           , S => n779, Z => n1298);
   U1749 : MUX2_X1 port map( A => n1298, B => n1297, S => n833, Z => n1299);
   U1750 : MUX2_X1 port map( A => n1299, B => n1296, S => n844, Z => n1300);
   U1751 : MUX2_X1 port map( A => n1300, B => n1293, S => n848, Z => n1301);
   U1752 : MUX2_X1 port map( A => REGISTERS_25_7_port, B => REGISTERS_26_7_port
                           , S => n779, Z => n1302);
   U1753 : MUX2_X1 port map( A => REGISTERS_23_7_port, B => REGISTERS_24_7_port
                           , S => n779, Z => n1303);
   U1754 : MUX2_X1 port map( A => n1303, B => n1302, S => n833, Z => n1304);
   U1755 : MUX2_X1 port map( A => REGISTERS_9_7_port, B => REGISTERS_10_7_port,
                           S => n779, Z => n1305);
   U1756 : MUX2_X1 port map( A => REGISTERS_7_7_port, B => REGISTERS_8_7_port, 
                           S => n785, Z => n1306);
   U1757 : MUX2_X1 port map( A => n1306, B => n1305, S => n834, Z => n1307);
   U1758 : MUX2_X1 port map( A => n1307, B => n1304, S => n844, Z => n1308);
   U1759 : MUX2_X1 port map( A => n1308, B => REGISTERS_39_7_port, S => n848, Z
                           => n1309);
   U1760 : MUX2_X1 port map( A => n1309, B => n1301, S => n302, Z => n1310);
   U1761 : MUX2_X1 port map( A => n1310, B => n1291, S => n301, Z => N12212);
   U1762 : MUX2_X1 port map( A => REGISTERS_5_8_port, B => REGISTERS_6_8_port, 
                           S => n803, Z => n1311);
   U1763 : MUX2_X1 port map( A => REGISTERS_3_8_port, B => REGISTERS_4_8_port, 
                           S => n804, Z => n1312);
   U1764 : MUX2_X1 port map( A => n1312, B => n1311, S => n834, Z => n1313);
   U1765 : MUX2_X1 port map( A => REGISTERS_37_8_port, B => REGISTERS_38_8_port
                           , S => n804, Z => n1314);
   U1766 : MUX2_X1 port map( A => REGISTERS_35_8_port, B => REGISTERS_36_8_port
                           , S => n804, Z => n1315);
   U1767 : MUX2_X1 port map( A => n1315, B => n1314, S => n834, Z => n1316);
   U1768 : MUX2_X1 port map( A => REGISTERS_21_8_port, B => REGISTERS_22_8_port
                           , S => n804, Z => n1317);
   U1769 : MUX2_X1 port map( A => REGISTERS_19_8_port, B => REGISTERS_20_8_port
                           , S => n804, Z => n1318);
   U1770 : MUX2_X1 port map( A => n1318, B => n1317, S => n834, Z => n1319);
   U1771 : MUX2_X1 port map( A => n1319, B => n1316, S => n844, Z => n1320);
   U1772 : MUX2_X1 port map( A => n1320, B => n1313, S => n848, Z => n1321);
   U1773 : MUX2_X1 port map( A => REGISTERS_29_8_port, B => REGISTERS_30_8_port
                           , S => n804, Z => n1322);
   U1774 : MUX2_X1 port map( A => REGISTERS_27_8_port, B => REGISTERS_28_8_port
                           , S => n804, Z => n1323);
   U1775 : MUX2_X1 port map( A => n1323, B => n1322, S => n834, Z => n1324);
   U1776 : MUX2_X1 port map( A => REGISTERS_13_8_port, B => REGISTERS_14_8_port
                           , S => n804, Z => n1325);
   U1777 : MUX2_X1 port map( A => REGISTERS_11_8_port, B => REGISTERS_12_8_port
                           , S => n804, Z => n1326);
   U1778 : MUX2_X1 port map( A => n1326, B => n1325, S => n834, Z => n1327);
   U1779 : MUX2_X1 port map( A => n1327, B => n1324, S => n844, Z => n1328);
   U1780 : MUX2_X1 port map( A => n1328, B => n1321, S => n302, Z => n1329);
   U1781 : MUX2_X1 port map( A => REGISTERS_1_8_port, B => REGISTERS_2_8_port, 
                           S => n803, Z => n1330);
   U1782 : MUX2_X1 port map( A => REGISTERS_0_8_port, B => n1330, S => n834, Z 
                           => n1331);
   U1783 : MUX2_X1 port map( A => REGISTERS_33_8_port, B => REGISTERS_34_8_port
                           , S => n803, Z => n1332);
   U1784 : MUX2_X1 port map( A => REGISTERS_31_8_port, B => REGISTERS_32_8_port
                           , S => n803, Z => n1333);
   U1785 : MUX2_X1 port map( A => n1333, B => n1332, S => n834, Z => n1334);
   U1786 : MUX2_X1 port map( A => REGISTERS_17_8_port, B => REGISTERS_18_8_port
                           , S => n803, Z => n1335);
   U1787 : MUX2_X1 port map( A => REGISTERS_15_8_port, B => REGISTERS_16_8_port
                           , S => n803, Z => n1336);
   U1788 : MUX2_X1 port map( A => n1336, B => n1335, S => n834, Z => n1337);
   U1789 : MUX2_X1 port map( A => n1337, B => n1334, S => n844, Z => n1338);
   U1790 : MUX2_X1 port map( A => n1338, B => n1331, S => n848, Z => n1339);
   U1791 : MUX2_X1 port map( A => REGISTERS_25_8_port, B => REGISTERS_26_8_port
                           , S => n802, Z => n1340);
   U1792 : MUX2_X1 port map( A => REGISTERS_23_8_port, B => REGISTERS_24_8_port
                           , S => n803, Z => n1341);
   U1793 : MUX2_X1 port map( A => n1341, B => n1340, S => n834, Z => n1342);
   U1794 : MUX2_X1 port map( A => REGISTERS_9_8_port, B => REGISTERS_10_8_port,
                           S => n803, Z => n1343);
   U1795 : MUX2_X1 port map( A => REGISTERS_7_8_port, B => REGISTERS_8_8_port, 
                           S => n803, Z => n1344);
   U1796 : MUX2_X1 port map( A => n1344, B => n1343, S => n834, Z => n1345);
   U1797 : MUX2_X1 port map( A => n1345, B => n1342, S => n844, Z => n1346);
   U1798 : MUX2_X1 port map( A => n1346, B => REGISTERS_39_8_port, S => n848, Z
                           => n1347);
   U1799 : MUX2_X1 port map( A => n1347, B => n1339, S => n302, Z => n1348);
   U1800 : MUX2_X1 port map( A => n1348, B => n1329, S => n301, Z => N12213);
   U1801 : MUX2_X1 port map( A => REGISTERS_5_9_port, B => REGISTERS_6_9_port, 
                           S => n803, Z => n1349);
   U1802 : MUX2_X1 port map( A => REGISTERS_3_9_port, B => REGISTERS_4_9_port, 
                           S => n803, Z => n1350);
   U1803 : MUX2_X1 port map( A => n1350, B => n1349, S => n835, Z => n1351);
   U1804 : MUX2_X1 port map( A => REGISTERS_37_9_port, B => REGISTERS_38_9_port
                           , S => n803, Z => n1352);
   U1805 : MUX2_X1 port map( A => REGISTERS_35_9_port, B => REGISTERS_36_9_port
                           , S => n802, Z => n1353);
   U1806 : MUX2_X1 port map( A => n1353, B => n1352, S => n835, Z => n1354);
   U1807 : MUX2_X1 port map( A => REGISTERS_21_9_port, B => REGISTERS_22_9_port
                           , S => n802, Z => n1355);
   U1808 : MUX2_X1 port map( A => REGISTERS_19_9_port, B => REGISTERS_20_9_port
                           , S => n802, Z => n1356);
   U1809 : MUX2_X1 port map( A => n1356, B => n1355, S => n835, Z => n1357);
   U1810 : MUX2_X1 port map( A => n1357, B => n1354, S => n844, Z => n1358);
   U1811 : MUX2_X1 port map( A => n1358, B => n1351, S => n848, Z => n1359);
   U1812 : MUX2_X1 port map( A => REGISTERS_29_9_port, B => REGISTERS_30_9_port
                           , S => n802, Z => n1360);
   U1813 : MUX2_X1 port map( A => REGISTERS_27_9_port, B => REGISTERS_28_9_port
                           , S => n802, Z => n1361);
   U1814 : MUX2_X1 port map( A => n1361, B => n1360, S => n835, Z => n1362);
   U1815 : MUX2_X1 port map( A => REGISTERS_13_9_port, B => REGISTERS_14_9_port
                           , S => n802, Z => n1363);
   U1816 : MUX2_X1 port map( A => REGISTERS_11_9_port, B => REGISTERS_12_9_port
                           , S => n802, Z => n1364);
   U1817 : MUX2_X1 port map( A => n1364, B => n1363, S => n835, Z => n1365);
   U1818 : MUX2_X1 port map( A => n1365, B => n1362, S => n844, Z => n1366);
   U1819 : MUX2_X1 port map( A => n1366, B => n1359, S => n302, Z => n1367);
   U1820 : MUX2_X1 port map( A => REGISTERS_1_9_port, B => REGISTERS_2_9_port, 
                           S => n802, Z => n1368);
   U1821 : MUX2_X1 port map( A => REGISTERS_0_9_port, B => n1368, S => n835, Z 
                           => n1369);
   U1822 : MUX2_X1 port map( A => REGISTERS_33_9_port, B => REGISTERS_34_9_port
                           , S => n801, Z => n1370);
   U1823 : MUX2_X1 port map( A => REGISTERS_31_9_port, B => REGISTERS_32_9_port
                           , S => n802, Z => n1371);
   U1824 : MUX2_X1 port map( A => n1371, B => n1370, S => n835, Z => n1372);
   U1825 : MUX2_X1 port map( A => REGISTERS_17_9_port, B => REGISTERS_18_9_port
                           , S => n802, Z => n1373);
   U1826 : MUX2_X1 port map( A => REGISTERS_15_9_port, B => REGISTERS_16_9_port
                           , S => n802, Z => n1374);
   U1827 : MUX2_X1 port map( A => n1374, B => n1373, S => n835, Z => n1375);
   U1828 : MUX2_X1 port map( A => n1375, B => n1372, S => n844, Z => n1376);
   U1829 : MUX2_X1 port map( A => n1376, B => n1369, S => n848, Z => n1377);
   U1830 : MUX2_X1 port map( A => REGISTERS_25_9_port, B => REGISTERS_26_9_port
                           , S => n801, Z => n1378);
   U1831 : MUX2_X1 port map( A => REGISTERS_23_9_port, B => REGISTERS_24_9_port
                           , S => n801, Z => n1379);
   U1832 : MUX2_X1 port map( A => n1379, B => n1378, S => n835, Z => n1380);
   U1833 : MUX2_X1 port map( A => REGISTERS_9_9_port, B => REGISTERS_10_9_port,
                           S => n801, Z => n1381);
   U1834 : MUX2_X1 port map( A => REGISTERS_7_9_port, B => REGISTERS_8_9_port, 
                           S => n801, Z => n1382);
   U1835 : MUX2_X1 port map( A => n1382, B => n1381, S => n835, Z => n1383);
   U1836 : MUX2_X1 port map( A => n1383, B => n1380, S => n844, Z => n1384);
   U1837 : MUX2_X1 port map( A => n1384, B => REGISTERS_39_9_port, S => n848, Z
                           => n1385);
   U1838 : MUX2_X1 port map( A => n1385, B => n1377, S => n302, Z => n1386);
   U1839 : MUX2_X1 port map( A => n1386, B => n1367, S => n301, Z => N12214);
   U1840 : MUX2_X1 port map( A => REGISTERS_5_10_port, B => REGISTERS_6_10_port
                           , S => n801, Z => n1387);
   U1841 : MUX2_X1 port map( A => REGISTERS_3_10_port, B => REGISTERS_4_10_port
                           , S => n801, Z => n1388);
   U1842 : MUX2_X1 port map( A => n1388, B => n1387, S => n835, Z => n1389);
   U1843 : MUX2_X1 port map( A => REGISTERS_37_10_port, B => 
                           REGISTERS_38_10_port, S => n801, Z => n1390);
   U1844 : MUX2_X1 port map( A => REGISTERS_35_10_port, B => 
                           REGISTERS_36_10_port, S => n801, Z => n1391);
   U1845 : MUX2_X1 port map( A => n1391, B => n1390, S => n835, Z => n1392);
   U1846 : MUX2_X1 port map( A => REGISTERS_21_10_port, B => 
                           REGISTERS_22_10_port, S => n801, Z => n1393);
   U1847 : MUX2_X1 port map( A => REGISTERS_19_10_port, B => 
                           REGISTERS_20_10_port, S => n801, Z => n1394);
   U1848 : MUX2_X1 port map( A => n1394, B => n1393, S => n836, Z => n1395);
   U1849 : MUX2_X1 port map( A => n1395, B => n1392, S => n844, Z => n1396);
   U1850 : MUX2_X1 port map( A => n1396, B => n1389, S => n848, Z => n1397);
   U1851 : MUX2_X1 port map( A => REGISTERS_29_10_port, B => 
                           REGISTERS_30_10_port, S => n801, Z => n1398);
   U1852 : MUX2_X1 port map( A => REGISTERS_27_10_port, B => 
                           REGISTERS_28_10_port, S => n799, Z => n1399);
   U1853 : MUX2_X1 port map( A => n1399, B => n1398, S => n836, Z => n1400);
   U1854 : MUX2_X1 port map( A => REGISTERS_13_10_port, B => 
                           REGISTERS_14_10_port, S => n800, Z => n1401);
   U1855 : MUX2_X1 port map( A => REGISTERS_11_10_port, B => 
                           REGISTERS_12_10_port, S => n800, Z => n1402);
   U1856 : MUX2_X1 port map( A => n1402, B => n1401, S => n836, Z => n1403);
   U1857 : MUX2_X1 port map( A => n1403, B => n1400, S => n844, Z => n1404);
   U1858 : MUX2_X1 port map( A => n1404, B => n1397, S => n302, Z => n1405);
   U1859 : MUX2_X1 port map( A => REGISTERS_1_10_port, B => REGISTERS_2_10_port
                           , S => n800, Z => n1406);
   U1860 : MUX2_X1 port map( A => REGISTERS_0_10_port, B => n1406, S => n836, Z
                           => n1407);
   U1861 : MUX2_X1 port map( A => REGISTERS_33_10_port, B => 
                           REGISTERS_34_10_port, S => n800, Z => n1408);
   U1862 : MUX2_X1 port map( A => REGISTERS_31_10_port, B => 
                           REGISTERS_32_10_port, S => n800, Z => n1409);
   U1863 : MUX2_X1 port map( A => n1409, B => n1408, S => n836, Z => n1410);
   U1864 : MUX2_X1 port map( A => REGISTERS_17_10_port, B => 
                           REGISTERS_18_10_port, S => n800, Z => n1411);
   U1865 : MUX2_X1 port map( A => REGISTERS_15_10_port, B => 
                           REGISTERS_16_10_port, S => n800, Z => n1412);
   U1866 : MUX2_X1 port map( A => n1412, B => n1411, S => n836, Z => n1413);
   U1867 : MUX2_X1 port map( A => n1413, B => n1410, S => n844, Z => n1414);
   U1868 : MUX2_X1 port map( A => n1414, B => n1407, S => n848, Z => n1415);
   U1869 : MUX2_X1 port map( A => REGISTERS_25_10_port, B => 
                           REGISTERS_26_10_port, S => n800, Z => n1416);
   U1870 : MUX2_X1 port map( A => REGISTERS_23_10_port, B => 
                           REGISTERS_24_10_port, S => n800, Z => n1417);
   U1871 : MUX2_X1 port map( A => n1417, B => n1416, S => n836, Z => n1418);
   U1872 : MUX2_X1 port map( A => REGISTERS_9_10_port, B => 
                           REGISTERS_10_10_port, S => n800, Z => n1419);
   U1873 : MUX2_X1 port map( A => REGISTERS_7_10_port, B => REGISTERS_8_10_port
                           , S => n800, Z => n1420);
   U1874 : MUX2_X1 port map( A => n1420, B => n1419, S => n836, Z => n1421);
   U1875 : MUX2_X1 port map( A => n1421, B => n1418, S => n844, Z => n1422);
   U1876 : MUX2_X1 port map( A => n1422, B => REGISTERS_39_10_port, S => n848, 
                           Z => n1423);
   U1877 : MUX2_X1 port map( A => n1423, B => n1415, S => n302, Z => n1424);
   U1878 : MUX2_X1 port map( A => n1424, B => n1405, S => n301, Z => N12215);
   U1879 : MUX2_X1 port map( A => REGISTERS_5_11_port, B => REGISTERS_6_11_port
                           , S => n800, Z => n1425);
   U1880 : MUX2_X1 port map( A => REGISTERS_3_11_port, B => REGISTERS_4_11_port
                           , S => n799, Z => n1426);
   U1881 : MUX2_X1 port map( A => n1426, B => n1425, S => n836, Z => n1427);
   U1882 : MUX2_X1 port map( A => REGISTERS_37_11_port, B => 
                           REGISTERS_38_11_port, S => n799, Z => n1428);
   U1883 : MUX2_X1 port map( A => REGISTERS_35_11_port, B => 
                           REGISTERS_36_11_port, S => n798, Z => n1429);
   U1884 : MUX2_X1 port map( A => n1429, B => n1428, S => n836, Z => n1430);
   U1885 : MUX2_X1 port map( A => REGISTERS_21_11_port, B => 
                           REGISTERS_22_11_port, S => n799, Z => n1431);
   U1886 : MUX2_X1 port map( A => REGISTERS_19_11_port, B => 
                           REGISTERS_20_11_port, S => n799, Z => n1432);
   U1887 : MUX2_X1 port map( A => n1432, B => n1431, S => n836, Z => n1433);
   U1888 : MUX2_X1 port map( A => n1433, B => n1430, S => n844, Z => n1434);
   U1889 : MUX2_X1 port map( A => n1434, B => n1427, S => n848, Z => n1435);
   U1890 : MUX2_X1 port map( A => REGISTERS_29_11_port, B => 
                           REGISTERS_30_11_port, S => n799, Z => n1436);
   U1891 : MUX2_X1 port map( A => REGISTERS_27_11_port, B => 
                           REGISTERS_28_11_port, S => n799, Z => n1437);
   U1892 : MUX2_X1 port map( A => n1437, B => n1436, S => n836, Z => n1438);
   U1893 : MUX2_X1 port map( A => REGISTERS_13_11_port, B => 
                           REGISTERS_14_11_port, S => n799, Z => n1439);
   U1894 : MUX2_X1 port map( A => REGISTERS_11_11_port, B => 
                           REGISTERS_12_11_port, S => n799, Z => n1440);
   U1895 : MUX2_X1 port map( A => n1440, B => n1439, S => n837, Z => n1441);
   U1896 : MUX2_X1 port map( A => n1441, B => n1438, S => n844, Z => n1442);
   U1897 : MUX2_X1 port map( A => n1442, B => n1435, S => n302, Z => n1443);
   U1898 : MUX2_X1 port map( A => REGISTERS_1_11_port, B => REGISTERS_2_11_port
                           , S => n799, Z => n1444);
   U1899 : MUX2_X1 port map( A => REGISTERS_0_11_port, B => n1444, S => n837, Z
                           => n1445);
   U1900 : MUX2_X1 port map( A => REGISTERS_33_11_port, B => 
                           REGISTERS_34_11_port, S => n799, Z => n1446);
   U1901 : MUX2_X1 port map( A => REGISTERS_31_11_port, B => 
                           REGISTERS_32_11_port, S => n799, Z => n1447);
   U1902 : MUX2_X1 port map( A => n1447, B => n1446, S => n837, Z => n1448);
   U1903 : MUX2_X1 port map( A => REGISTERS_17_11_port, B => 
                           REGISTERS_18_11_port, S => n798, Z => n1449);
   U1904 : MUX2_X1 port map( A => REGISTERS_15_11_port, B => 
                           REGISTERS_16_11_port, S => n798, Z => n1450);
   U1905 : MUX2_X1 port map( A => n1450, B => n1449, S => n837, Z => n1451);
   U1906 : MUX2_X1 port map( A => n1451, B => n1448, S => n844, Z => n1452);
   U1907 : MUX2_X1 port map( A => n1452, B => n1445, S => n848, Z => n1453);
   U1908 : MUX2_X1 port map( A => REGISTERS_25_11_port, B => 
                           REGISTERS_26_11_port, S => n798, Z => n1454);
   U1909 : MUX2_X1 port map( A => REGISTERS_23_11_port, B => 
                           REGISTERS_24_11_port, S => n798, Z => n1455);
   U1910 : MUX2_X1 port map( A => n1455, B => n1454, S => n837, Z => n1456);
   U1911 : MUX2_X1 port map( A => REGISTERS_9_11_port, B => 
                           REGISTERS_10_11_port, S => n798, Z => n1457);
   U1912 : MUX2_X1 port map( A => REGISTERS_7_11_port, B => REGISTERS_8_11_port
                           , S => n798, Z => n1458);
   U1913 : MUX2_X1 port map( A => n1458, B => n1457, S => n837, Z => n1459);
   U1914 : MUX2_X1 port map( A => n1459, B => n1456, S => n844, Z => n1460);
   U1915 : MUX2_X1 port map( A => n1460, B => REGISTERS_39_11_port, S => n848, 
                           Z => n1461);
   U1916 : MUX2_X1 port map( A => n1461, B => n1453, S => n302, Z => n1462);
   U1917 : MUX2_X1 port map( A => n1462, B => n1443, S => n301, Z => N12216);
   U1918 : MUX2_X1 port map( A => REGISTERS_5_12_port, B => REGISTERS_6_12_port
                           , S => n798, Z => n1463);
   U1919 : MUX2_X1 port map( A => REGISTERS_3_12_port, B => REGISTERS_4_12_port
                           , S => n798, Z => n1464);
   U1920 : MUX2_X1 port map( A => n1464, B => n1463, S => n837, Z => n1465);
   U1921 : MUX2_X1 port map( A => REGISTERS_37_12_port, B => 
                           REGISTERS_38_12_port, S => n798, Z => n1466);
   U1922 : MUX2_X1 port map( A => REGISTERS_35_12_port, B => 
                           REGISTERS_36_12_port, S => n798, Z => n1467);
   U1923 : MUX2_X1 port map( A => n1467, B => n1466, S => n837, Z => n1468);
   U1924 : MUX2_X1 port map( A => REGISTERS_21_12_port, B => 
                           REGISTERS_22_12_port, S => n797, Z => n1469);
   U1925 : MUX2_X1 port map( A => REGISTERS_19_12_port, B => 
                           REGISTERS_20_12_port, S => n797, Z => n1470);
   U1926 : MUX2_X1 port map( A => n1470, B => n1469, S => n837, Z => n1471);
   U1927 : MUX2_X1 port map( A => n1471, B => n1468, S => n844, Z => n1472);
   U1928 : MUX2_X1 port map( A => n1472, B => n1465, S => n848, Z => n1473);
   U1929 : MUX2_X1 port map( A => REGISTERS_29_12_port, B => 
                           REGISTERS_30_12_port, S => n797, Z => n1474);
   U1930 : MUX2_X1 port map( A => REGISTERS_27_12_port, B => 
                           REGISTERS_28_12_port, S => n797, Z => n1475);
   U1931 : MUX2_X1 port map( A => n1475, B => n1474, S => n837, Z => n1476);
   U1932 : MUX2_X1 port map( A => REGISTERS_13_12_port, B => 
                           REGISTERS_14_12_port, S => n797, Z => n1477);
   U1933 : MUX2_X1 port map( A => REGISTERS_11_12_port, B => 
                           REGISTERS_12_12_port, S => n797, Z => n1478);
   U1934 : MUX2_X1 port map( A => n1478, B => n1477, S => n837, Z => n1479);
   U1935 : MUX2_X1 port map( A => n1479, B => n1476, S => n844, Z => n1480);
   U1936 : MUX2_X1 port map( A => n1480, B => n1473, S => n302, Z => n1481);
   U1937 : MUX2_X1 port map( A => REGISTERS_1_12_port, B => REGISTERS_2_12_port
                           , S => n797, Z => n1482);
   U1938 : MUX2_X1 port map( A => REGISTERS_0_12_port, B => n1482, S => n837, Z
                           => n1483);
   U1939 : MUX2_X1 port map( A => REGISTERS_33_12_port, B => 
                           REGISTERS_34_12_port, S => n797, Z => n1484);
   U1940 : MUX2_X1 port map( A => REGISTERS_31_12_port, B => 
                           REGISTERS_32_12_port, S => n797, Z => n1485);
   U1941 : MUX2_X1 port map( A => n1485, B => n1484, S => n838, Z => n1486);
   U1942 : MUX2_X1 port map( A => REGISTERS_17_12_port, B => 
                           REGISTERS_18_12_port, S => n797, Z => n1487);
   U1943 : MUX2_X1 port map( A => REGISTERS_15_12_port, B => 
                           REGISTERS_16_12_port, S => n797, Z => n1488);
   U1944 : MUX2_X1 port map( A => n1488, B => n1487, S => n838, Z => n1489);
   U1945 : MUX2_X1 port map( A => n1489, B => n1486, S => n844, Z => n1490);
   U1946 : MUX2_X1 port map( A => n1490, B => n1483, S => n848, Z => n1491);
   U1947 : MUX2_X1 port map( A => REGISTERS_25_12_port, B => 
                           REGISTERS_26_12_port, S => n797, Z => n1492);
   U1948 : MUX2_X1 port map( A => REGISTERS_23_12_port, B => 
                           REGISTERS_24_12_port, S => n796, Z => n1493);
   U1949 : MUX2_X1 port map( A => n1493, B => n1492, S => n838, Z => n1494);
   U1950 : MUX2_X1 port map( A => REGISTERS_9_12_port, B => 
                           REGISTERS_10_12_port, S => n796, Z => n1495);
   U1951 : MUX2_X1 port map( A => REGISTERS_7_12_port, B => REGISTERS_8_12_port
                           , S => n796, Z => n1496);
   U1952 : MUX2_X1 port map( A => n1496, B => n1495, S => n838, Z => n1497);
   U1953 : MUX2_X1 port map( A => n1497, B => n1494, S => n844, Z => n1498);
   U1954 : MUX2_X1 port map( A => n1498, B => REGISTERS_39_12_port, S => n848, 
                           Z => n1499);
   U1955 : MUX2_X1 port map( A => n1499, B => n1491, S => n302, Z => n1500);
   U1956 : MUX2_X1 port map( A => n1500, B => n1481, S => n301, Z => N12217);
   U1957 : MUX2_X1 port map( A => REGISTERS_5_13_port, B => REGISTERS_6_13_port
                           , S => n796, Z => n1501);
   U1958 : MUX2_X1 port map( A => REGISTERS_3_13_port, B => REGISTERS_4_13_port
                           , S => n796, Z => n1502);
   U1959 : MUX2_X1 port map( A => n1502, B => n1501, S => n838, Z => n1503);
   U1960 : MUX2_X1 port map( A => REGISTERS_37_13_port, B => 
                           REGISTERS_38_13_port, S => n796, Z => n1504);
   U1961 : MUX2_X1 port map( A => REGISTERS_35_13_port, B => 
                           REGISTERS_36_13_port, S => n796, Z => n1505);
   U1962 : MUX2_X1 port map( A => n1505, B => n1504, S => n838, Z => n1506);
   U1963 : MUX2_X1 port map( A => REGISTERS_21_13_port, B => 
                           REGISTERS_22_13_port, S => n796, Z => n1507);
   U1964 : MUX2_X1 port map( A => REGISTERS_19_13_port, B => 
                           REGISTERS_20_13_port, S => n796, Z => n1508);
   U1965 : MUX2_X1 port map( A => n1508, B => n1507, S => n838, Z => n1509);
   U1966 : MUX2_X1 port map( A => n1509, B => n1506, S => n844, Z => n1510);
   U1967 : MUX2_X1 port map( A => n1510, B => n1503, S => n848, Z => n1511);
   U1968 : MUX2_X1 port map( A => REGISTERS_29_13_port, B => 
                           REGISTERS_30_13_port, S => n796, Z => n1512);
   U1969 : MUX2_X1 port map( A => REGISTERS_27_13_port, B => 
                           REGISTERS_28_13_port, S => n796, Z => n1513);
   U1970 : MUX2_X1 port map( A => n1513, B => n1512, S => n838, Z => n1514);
   U1971 : MUX2_X1 port map( A => REGISTERS_13_13_port, B => 
                           REGISTERS_14_13_port, S => n796, Z => n1515);
   U1972 : MUX2_X1 port map( A => REGISTERS_11_13_port, B => 
                           REGISTERS_12_13_port, S => n795, Z => n1516);
   U1973 : MUX2_X1 port map( A => n1516, B => n1515, S => n838, Z => n1517);
   U1974 : MUX2_X1 port map( A => n1517, B => n1514, S => n844, Z => n1518);
   U1975 : MUX2_X1 port map( A => n1518, B => n1511, S => n302, Z => n1519);
   U1976 : MUX2_X1 port map( A => REGISTERS_1_13_port, B => REGISTERS_2_13_port
                           , S => n795, Z => n1520);
   U1977 : MUX2_X1 port map( A => REGISTERS_0_13_port, B => n1520, S => n838, Z
                           => n1521);
   U1978 : MUX2_X1 port map( A => REGISTERS_33_13_port, B => 
                           REGISTERS_34_13_port, S => n795, Z => n1522);
   U1979 : MUX2_X1 port map( A => REGISTERS_31_13_port, B => 
                           REGISTERS_32_13_port, S => n795, Z => n1523);
   U1980 : MUX2_X1 port map( A => n1523, B => n1522, S => n838, Z => n1524);
   U1981 : MUX2_X1 port map( A => REGISTERS_17_13_port, B => 
                           REGISTERS_18_13_port, S => n795, Z => n1525);
   U1982 : MUX2_X1 port map( A => REGISTERS_15_13_port, B => 
                           REGISTERS_16_13_port, S => n795, Z => n1526);
   U1983 : MUX2_X1 port map( A => n1526, B => n1525, S => n838, Z => n1527);
   U1984 : MUX2_X1 port map( A => n1527, B => n1524, S => n843, Z => n1528);
   U1985 : MUX2_X1 port map( A => n1528, B => n1521, S => n848, Z => n1529);
   U1986 : MUX2_X1 port map( A => REGISTERS_25_13_port, B => 
                           REGISTERS_26_13_port, S => n795, Z => n1530);
   U1987 : MUX2_X1 port map( A => REGISTERS_23_13_port, B => 
                           REGISTERS_24_13_port, S => n795, Z => n1531);
   U1988 : MUX2_X1 port map( A => n1531, B => n1530, S => n839, Z => n1532);
   U1989 : MUX2_X1 port map( A => REGISTERS_9_13_port, B => 
                           REGISTERS_10_13_port, S => n795, Z => n1533);
   U1990 : MUX2_X1 port map( A => REGISTERS_7_13_port, B => REGISTERS_8_13_port
                           , S => n795, Z => n1534);
   U1991 : MUX2_X1 port map( A => n1534, B => n1533, S => n839, Z => n1535);
   U1992 : MUX2_X1 port map( A => n1535, B => n1532, S => n843, Z => n1536);
   U1993 : MUX2_X1 port map( A => n1536, B => REGISTERS_39_13_port, S => n848, 
                           Z => n1537);
   U1994 : MUX2_X1 port map( A => n1537, B => n1529, S => n302, Z => n1538);
   U1995 : MUX2_X1 port map( A => n1538, B => n1519, S => n301, Z => N12218);
   U1996 : MUX2_X1 port map( A => REGISTERS_5_14_port, B => REGISTERS_6_14_port
                           , S => n795, Z => n1539);
   U1997 : MUX2_X1 port map( A => REGISTERS_3_14_port, B => REGISTERS_4_14_port
                           , S => n795, Z => n1540);
   U1998 : MUX2_X1 port map( A => n1540, B => n1539, S => n839, Z => n1541);
   U1999 : MUX2_X1 port map( A => REGISTERS_37_14_port, B => 
                           REGISTERS_38_14_port, S => n794, Z => n1542);
   U2000 : MUX2_X1 port map( A => REGISTERS_35_14_port, B => 
                           REGISTERS_36_14_port, S => n794, Z => n1543);
   U2001 : MUX2_X1 port map( A => n1543, B => n1542, S => n839, Z => n1544);
   U2002 : MUX2_X1 port map( A => REGISTERS_21_14_port, B => 
                           REGISTERS_22_14_port, S => n794, Z => n1545);
   U2003 : MUX2_X1 port map( A => REGISTERS_19_14_port, B => 
                           REGISTERS_20_14_port, S => n794, Z => n1546);
   U2004 : MUX2_X1 port map( A => n1546, B => n1545, S => n839, Z => n1547);
   U2005 : MUX2_X1 port map( A => n1547, B => n1544, S => n843, Z => n1548);
   U2006 : MUX2_X1 port map( A => n1548, B => n1541, S => n848, Z => n1549);
   U2007 : MUX2_X1 port map( A => REGISTERS_29_14_port, B => 
                           REGISTERS_30_14_port, S => n794, Z => n1550);
   U2008 : MUX2_X1 port map( A => REGISTERS_27_14_port, B => 
                           REGISTERS_28_14_port, S => n794, Z => n1551);
   U2009 : MUX2_X1 port map( A => n1551, B => n1550, S => n839, Z => n1552);
   U2010 : MUX2_X1 port map( A => REGISTERS_13_14_port, B => 
                           REGISTERS_14_14_port, S => n794, Z => n1553);
   U2011 : MUX2_X1 port map( A => REGISTERS_11_14_port, B => 
                           REGISTERS_12_14_port, S => n794, Z => n1554);
   U2012 : MUX2_X1 port map( A => n1554, B => n1553, S => n839, Z => n1555);
   U2013 : MUX2_X1 port map( A => n1555, B => n1552, S => n843, Z => n1556);
   U2014 : MUX2_X1 port map( A => n1556, B => n1549, S => n302, Z => n1557);
   U2015 : MUX2_X1 port map( A => REGISTERS_1_14_port, B => REGISTERS_2_14_port
                           , S => n794, Z => n1558);
   U2016 : MUX2_X1 port map( A => REGISTERS_0_14_port, B => n1558, S => n839, Z
                           => n1559);
   U2017 : MUX2_X1 port map( A => REGISTERS_33_14_port, B => 
                           REGISTERS_34_14_port, S => n794, Z => n1560);
   U2018 : MUX2_X1 port map( A => REGISTERS_31_14_port, B => 
                           REGISTERS_32_14_port, S => n794, Z => n1561);
   U2019 : MUX2_X1 port map( A => n1561, B => n1560, S => n839, Z => n1562);
   U2020 : MUX2_X1 port map( A => REGISTERS_17_14_port, B => 
                           REGISTERS_18_14_port, S => n794, Z => n1563);
   U2021 : MUX2_X1 port map( A => REGISTERS_15_14_port, B => 
                           REGISTERS_16_14_port, S => n793, Z => n1564);
   U2022 : MUX2_X1 port map( A => n1564, B => n1563, S => n839, Z => n1565);
   U2023 : MUX2_X1 port map( A => n1565, B => n1562, S => n843, Z => n1566);
   U2024 : MUX2_X1 port map( A => n1566, B => n1559, S => n848, Z => n1567);
   U2025 : MUX2_X1 port map( A => REGISTERS_25_14_port, B => 
                           REGISTERS_26_14_port, S => n793, Z => n1568);
   U2026 : MUX2_X1 port map( A => REGISTERS_23_14_port, B => 
                           REGISTERS_24_14_port, S => n793, Z => n1569);
   U2027 : MUX2_X1 port map( A => n1569, B => n1568, S => n839, Z => n1570);
   U2028 : MUX2_X1 port map( A => REGISTERS_9_14_port, B => 
                           REGISTERS_10_14_port, S => n793, Z => n1571);
   U2029 : MUX2_X1 port map( A => REGISTERS_7_14_port, B => REGISTERS_8_14_port
                           , S => n793, Z => n1572);
   U2030 : MUX2_X1 port map( A => n1572, B => n1571, S => n839, Z => n1573);
   U2031 : MUX2_X1 port map( A => n1573, B => n1570, S => n843, Z => n1574);
   U2032 : MUX2_X1 port map( A => n1574, B => REGISTERS_39_14_port, S => n848, 
                           Z => n1575);
   U2033 : MUX2_X1 port map( A => n1575, B => n1567, S => n302, Z => n1576);
   U2034 : MUX2_X1 port map( A => n1576, B => n1557, S => n301, Z => N12219);
   U2035 : MUX2_X1 port map( A => REGISTERS_5_15_port, B => REGISTERS_6_15_port
                           , S => n793, Z => n1577);
   U2036 : MUX2_X1 port map( A => REGISTERS_3_15_port, B => REGISTERS_4_15_port
                           , S => n793, Z => n1578);
   U2037 : MUX2_X1 port map( A => n1578, B => n1577, S => n840, Z => n1579);
   U2038 : MUX2_X1 port map( A => REGISTERS_37_15_port, B => 
                           REGISTERS_38_15_port, S => n793, Z => n1580);
   U2039 : MUX2_X1 port map( A => REGISTERS_35_15_port, B => 
                           REGISTERS_36_15_port, S => n793, Z => n1581);
   U2040 : MUX2_X1 port map( A => n1581, B => n1580, S => n840, Z => n1582);
   U2041 : MUX2_X1 port map( A => REGISTERS_21_15_port, B => 
                           REGISTERS_22_15_port, S => n793, Z => n1583);
   U2042 : MUX2_X1 port map( A => REGISTERS_19_15_port, B => 
                           REGISTERS_20_15_port, S => n793, Z => n1584);
   U2043 : MUX2_X1 port map( A => n1584, B => n1583, S => n840, Z => n1585);
   U2044 : MUX2_X1 port map( A => n1585, B => n1582, S => n843, Z => n1586);
   U2045 : MUX2_X1 port map( A => n1586, B => n1579, S => n848, Z => n1587);
   U2046 : MUX2_X1 port map( A => REGISTERS_29_15_port, B => 
                           REGISTERS_30_15_port, S => n793, Z => n1588);
   U2047 : MUX2_X1 port map( A => REGISTERS_27_15_port, B => 
                           REGISTERS_28_15_port, S => n792, Z => n1589);
   U2048 : MUX2_X1 port map( A => n1589, B => n1588, S => n840, Z => n1590);
   U2049 : MUX2_X1 port map( A => REGISTERS_13_15_port, B => 
                           REGISTERS_14_15_port, S => n792, Z => n1591);
   U2050 : MUX2_X1 port map( A => REGISTERS_11_15_port, B => 
                           REGISTERS_12_15_port, S => n792, Z => n1592);
   U2051 : MUX2_X1 port map( A => n1592, B => n1591, S => n840, Z => n1593);
   U2052 : MUX2_X1 port map( A => n1593, B => n1590, S => n843, Z => n1594);
   U2053 : MUX2_X1 port map( A => n1594, B => n1587, S => n302, Z => n1595);
   U2054 : MUX2_X1 port map( A => REGISTERS_1_15_port, B => REGISTERS_2_15_port
                           , S => n792, Z => n1596);
   U2055 : MUX2_X1 port map( A => REGISTERS_0_15_port, B => n1596, S => n840, Z
                           => n1597);
   U2056 : MUX2_X1 port map( A => REGISTERS_33_15_port, B => 
                           REGISTERS_34_15_port, S => n792, Z => n1598);
   U2057 : MUX2_X1 port map( A => REGISTERS_31_15_port, B => 
                           REGISTERS_32_15_port, S => n792, Z => n1599);
   U2058 : MUX2_X1 port map( A => n1599, B => n1598, S => n840, Z => n1600);
   U2059 : MUX2_X1 port map( A => REGISTERS_17_15_port, B => 
                           REGISTERS_18_15_port, S => n792, Z => n1601);
   U2060 : MUX2_X1 port map( A => REGISTERS_15_15_port, B => 
                           REGISTERS_16_15_port, S => n792, Z => n1602);
   U2061 : MUX2_X1 port map( A => n1602, B => n1601, S => n840, Z => n1603);
   U2062 : MUX2_X1 port map( A => n1603, B => n1600, S => n843, Z => n1604);
   U2063 : MUX2_X1 port map( A => n1604, B => n1597, S => n848, Z => n1605);
   U2064 : MUX2_X1 port map( A => REGISTERS_25_15_port, B => 
                           REGISTERS_26_15_port, S => n792, Z => n1606);
   U2065 : MUX2_X1 port map( A => REGISTERS_23_15_port, B => 
                           REGISTERS_24_15_port, S => n792, Z => n1607);
   U2066 : MUX2_X1 port map( A => n1607, B => n1606, S => n840, Z => n1608);
   U2067 : MUX2_X1 port map( A => REGISTERS_9_15_port, B => 
                           REGISTERS_10_15_port, S => n798, Z => n1609);
   U2068 : MUX2_X1 port map( A => REGISTERS_7_15_port, B => REGISTERS_8_15_port
                           , S => n766, Z => n1610);
   U2069 : MUX2_X1 port map( A => n1610, B => n1609, S => n820, Z => n1611);
   U2070 : MUX2_X1 port map( A => n1611, B => n1608, S => n843, Z => n1612);
   U2071 : MUX2_X1 port map( A => n1612, B => REGISTERS_39_15_port, S => n848, 
                           Z => n1613);
   U2072 : MUX2_X1 port map( A => n1613, B => n1605, S => n302, Z => n1614);
   U2073 : MUX2_X1 port map( A => n1614, B => n1595, S => n301, Z => N12220);
   U2074 : MUX2_X1 port map( A => REGISTERS_5_16_port, B => REGISTERS_6_16_port
                           , S => n766, Z => n1615);
   U2075 : MUX2_X1 port map( A => REGISTERS_3_16_port, B => REGISTERS_4_16_port
                           , S => n766, Z => n1616);
   U2076 : MUX2_X1 port map( A => n1616, B => n1615, S => n814, Z => n1617);
   U2077 : MUX2_X1 port map( A => REGISTERS_37_16_port, B => 
                           REGISTERS_38_16_port, S => n766, Z => n1618);
   U2078 : MUX2_X1 port map( A => REGISTERS_35_16_port, B => 
                           REGISTERS_36_16_port, S => n766, Z => n1619);
   U2079 : MUX2_X1 port map( A => n1619, B => n1618, S => n814, Z => n1620);
   U2080 : MUX2_X1 port map( A => REGISTERS_21_16_port, B => 
                           REGISTERS_22_16_port, S => n766, Z => n1621);
   U2081 : MUX2_X1 port map( A => REGISTERS_19_16_port, B => 
                           REGISTERS_20_16_port, S => n766, Z => n1622);
   U2082 : MUX2_X1 port map( A => n1622, B => n1621, S => n814, Z => n1623);
   U2083 : MUX2_X1 port map( A => n1623, B => n1620, S => n843, Z => n1624);
   U2084 : MUX2_X1 port map( A => n1624, B => n1617, S => n848, Z => n1625);
   U2085 : MUX2_X1 port map( A => REGISTERS_29_16_port, B => 
                           REGISTERS_30_16_port, S => n766, Z => n1626);
   U2086 : MUX2_X1 port map( A => REGISTERS_27_16_port, B => 
                           REGISTERS_28_16_port, S => n766, Z => n1627);
   U2087 : MUX2_X1 port map( A => n1627, B => n1626, S => n814, Z => n1628);
   U2088 : MUX2_X1 port map( A => REGISTERS_13_16_port, B => 
                           REGISTERS_14_16_port, S => n766, Z => n1629);
   U2089 : MUX2_X1 port map( A => REGISTERS_11_16_port, B => 
                           REGISTERS_12_16_port, S => n765, Z => n1630);
   U2090 : MUX2_X1 port map( A => n1630, B => n1629, S => n814, Z => n1631);
   U2091 : MUX2_X1 port map( A => n1631, B => n1628, S => n843, Z => n1632);
   U2092 : MUX2_X1 port map( A => n1632, B => n1625, S => n302, Z => n1633);
   U2093 : MUX2_X1 port map( A => REGISTERS_1_16_port, B => REGISTERS_2_16_port
                           , S => n765, Z => n1634);
   U2094 : MUX2_X1 port map( A => REGISTERS_0_16_port, B => n1634, S => n814, Z
                           => n1635);
   U2095 : MUX2_X1 port map( A => REGISTERS_33_16_port, B => 
                           REGISTERS_34_16_port, S => n765, Z => n1636);
   U2096 : MUX2_X1 port map( A => REGISTERS_31_16_port, B => 
                           REGISTERS_32_16_port, S => n765, Z => n1637);
   U2097 : MUX2_X1 port map( A => n1637, B => n1636, S => n814, Z => n1638);
   U2098 : MUX2_X1 port map( A => REGISTERS_17_16_port, B => 
                           REGISTERS_18_16_port, S => n765, Z => n1639);
   U2099 : MUX2_X1 port map( A => REGISTERS_15_16_port, B => 
                           REGISTERS_16_16_port, S => n765, Z => n1640);
   U2100 : MUX2_X1 port map( A => n1640, B => n1639, S => n814, Z => n1641);
   U2101 : MUX2_X1 port map( A => n1641, B => n1638, S => n843, Z => n1642);
   U2102 : MUX2_X1 port map( A => n1642, B => n1635, S => n848, Z => n1643);
   U2103 : MUX2_X1 port map( A => REGISTERS_25_16_port, B => 
                           REGISTERS_26_16_port, S => n765, Z => n1644);
   U2104 : MUX2_X1 port map( A => REGISTERS_23_16_port, B => 
                           REGISTERS_24_16_port, S => n765, Z => n1645);
   U2105 : MUX2_X1 port map( A => n1645, B => n1644, S => n814, Z => n1646);
   U2106 : MUX2_X1 port map( A => REGISTERS_9_16_port, B => 
                           REGISTERS_10_16_port, S => n765, Z => n1647);
   U2107 : MUX2_X1 port map( A => REGISTERS_7_16_port, B => REGISTERS_8_16_port
                           , S => n765, Z => n1648);
   U2108 : MUX2_X1 port map( A => n1648, B => n1647, S => n814, Z => n1649);
   U2109 : MUX2_X1 port map( A => n1649, B => n1646, S => n843, Z => n1650);
   U2110 : MUX2_X1 port map( A => n1650, B => REGISTERS_39_16_port, S => n848, 
                           Z => n1651);
   U2111 : MUX2_X1 port map( A => n1651, B => n1643, S => n302, Z => n1652);
   U2112 : MUX2_X1 port map( A => n1652, B => n1633, S => n301, Z => N12221);
   U2113 : MUX2_X1 port map( A => REGISTERS_5_17_port, B => REGISTERS_6_17_port
                           , S => n765, Z => n1653);
   U2114 : MUX2_X1 port map( A => REGISTERS_3_17_port, B => REGISTERS_4_17_port
                           , S => n765, Z => n1654);
   U2115 : MUX2_X1 port map( A => n1654, B => n1653, S => n815, Z => n1655);
   U2116 : MUX2_X1 port map( A => REGISTERS_37_17_port, B => 
                           REGISTERS_38_17_port, S => n764, Z => n1656);
   U2117 : MUX2_X1 port map( A => REGISTERS_35_17_port, B => 
                           REGISTERS_36_17_port, S => n764, Z => n1657);
   U2118 : MUX2_X1 port map( A => n1657, B => n1656, S => n815, Z => n1658);
   U2119 : MUX2_X1 port map( A => REGISTERS_21_17_port, B => 
                           REGISTERS_22_17_port, S => n764, Z => n1659);
   U2120 : MUX2_X1 port map( A => REGISTERS_19_17_port, B => 
                           REGISTERS_20_17_port, S => n764, Z => n1660);
   U2121 : MUX2_X1 port map( A => n1660, B => n1659, S => n815, Z => n1661);
   U2122 : MUX2_X1 port map( A => n1661, B => n1658, S => n843, Z => n1662);
   U2123 : MUX2_X1 port map( A => n1662, B => n1655, S => n848, Z => n1663);
   U2124 : MUX2_X1 port map( A => REGISTERS_29_17_port, B => 
                           REGISTERS_30_17_port, S => n764, Z => n1664);
   U2125 : MUX2_X1 port map( A => REGISTERS_27_17_port, B => 
                           REGISTERS_28_17_port, S => n764, Z => n1665);
   U2126 : MUX2_X1 port map( A => n1665, B => n1664, S => n815, Z => n1666);
   U2127 : MUX2_X1 port map( A => REGISTERS_13_17_port, B => 
                           REGISTERS_14_17_port, S => n764, Z => n1667);
   U2128 : MUX2_X1 port map( A => REGISTERS_11_17_port, B => 
                           REGISTERS_12_17_port, S => n764, Z => n1668);
   U2129 : MUX2_X1 port map( A => n1668, B => n1667, S => n815, Z => n1669);
   U2130 : MUX2_X1 port map( A => n1669, B => n1666, S => n843, Z => n1670);
   U2131 : MUX2_X1 port map( A => n1670, B => n1663, S => n302, Z => n1671);
   U2132 : MUX2_X1 port map( A => REGISTERS_1_17_port, B => REGISTERS_2_17_port
                           , S => n764, Z => n1672);
   U2133 : MUX2_X1 port map( A => REGISTERS_0_17_port, B => n1672, S => n815, Z
                           => n1673);
   U2134 : MUX2_X1 port map( A => REGISTERS_33_17_port, B => 
                           REGISTERS_34_17_port, S => n764, Z => n1674);
   U2135 : MUX2_X1 port map( A => REGISTERS_31_17_port, B => 
                           REGISTERS_32_17_port, S => n764, Z => n1675);
   U2136 : MUX2_X1 port map( A => n1675, B => n1674, S => n815, Z => n1676);
   U2137 : MUX2_X1 port map( A => REGISTERS_17_17_port, B => 
                           REGISTERS_18_17_port, S => n764, Z => n1677);
   U2138 : MUX2_X1 port map( A => REGISTERS_15_17_port, B => 
                           REGISTERS_16_17_port, S => n763, Z => n1678);
   U2139 : MUX2_X1 port map( A => n1678, B => n1677, S => n815, Z => n1679);
   U2140 : MUX2_X1 port map( A => n1679, B => n1676, S => n843, Z => n1680);
   U2141 : MUX2_X1 port map( A => n1680, B => n1673, S => n848, Z => n1681);
   U2142 : MUX2_X1 port map( A => REGISTERS_25_17_port, B => 
                           REGISTERS_26_17_port, S => n763, Z => n1682);
   U2143 : MUX2_X1 port map( A => REGISTERS_23_17_port, B => 
                           REGISTERS_24_17_port, S => n763, Z => n1683);
   U2144 : MUX2_X1 port map( A => n1683, B => n1682, S => n815, Z => n1684);
   U2145 : MUX2_X1 port map( A => REGISTERS_9_17_port, B => 
                           REGISTERS_10_17_port, S => n763, Z => n1685);
   U2146 : MUX2_X1 port map( A => REGISTERS_7_17_port, B => REGISTERS_8_17_port
                           , S => n763, Z => n1686);
   U2147 : MUX2_X1 port map( A => n1686, B => n1685, S => n815, Z => n1687);
   U2148 : MUX2_X1 port map( A => n1687, B => n1684, S => n843, Z => n1688);
   U2149 : MUX2_X1 port map( A => n1688, B => REGISTERS_39_17_port, S => n848, 
                           Z => n1689);
   U2150 : MUX2_X1 port map( A => n1689, B => n1681, S => n302, Z => n1690);
   U2151 : MUX2_X1 port map( A => n1690, B => n1671, S => n301, Z => N12222);
   U2152 : MUX2_X1 port map( A => REGISTERS_5_18_port, B => REGISTERS_6_18_port
                           , S => n763, Z => n1691);
   U2153 : MUX2_X1 port map( A => REGISTERS_3_18_port, B => REGISTERS_4_18_port
                           , S => n763, Z => n1692);
   U2154 : MUX2_X1 port map( A => n1692, B => n1691, S => n815, Z => n1693);
   U2155 : MUX2_X1 port map( A => REGISTERS_37_18_port, B => 
                           REGISTERS_38_18_port, S => n763, Z => n1694);
   U2156 : MUX2_X1 port map( A => REGISTERS_35_18_port, B => 
                           REGISTERS_36_18_port, S => n763, Z => n1695);
   U2157 : MUX2_X1 port map( A => n1695, B => n1694, S => n815, Z => n1696);
   U2158 : MUX2_X1 port map( A => REGISTERS_21_18_port, B => 
                           REGISTERS_22_18_port, S => n763, Z => n1697);
   U2159 : MUX2_X1 port map( A => REGISTERS_19_18_port, B => 
                           REGISTERS_20_18_port, S => n763, Z => n1698);
   U2160 : MUX2_X1 port map( A => n1698, B => n1697, S => n816, Z => n1699);
   U2161 : MUX2_X1 port map( A => n1699, B => n1696, S => n843, Z => n1700);
   U2162 : MUX2_X1 port map( A => n1700, B => n1693, S => n848, Z => n1701);
   U2163 : MUX2_X1 port map( A => REGISTERS_29_18_port, B => 
                           REGISTERS_30_18_port, S => n763, Z => n1702);
   U2164 : MUX2_X1 port map( A => REGISTERS_27_18_port, B => 
                           REGISTERS_28_18_port, S => n762, Z => n1703);
   U2165 : MUX2_X1 port map( A => n1703, B => n1702, S => n816, Z => n1704);
   U2166 : MUX2_X1 port map( A => REGISTERS_13_18_port, B => 
                           REGISTERS_14_18_port, S => n762, Z => n1705);
   U2167 : MUX2_X1 port map( A => REGISTERS_11_18_port, B => 
                           REGISTERS_12_18_port, S => n762, Z => n1706);
   U2168 : MUX2_X1 port map( A => n1706, B => n1705, S => n816, Z => n1707);
   U2169 : MUX2_X1 port map( A => n1707, B => n1704, S => n843, Z => n1708);
   U2170 : MUX2_X1 port map( A => n1708, B => n1701, S => n302, Z => n1709);
   U2171 : MUX2_X1 port map( A => REGISTERS_1_18_port, B => REGISTERS_2_18_port
                           , S => n762, Z => n1710);
   U2172 : MUX2_X1 port map( A => REGISTERS_0_18_port, B => n1710, S => n816, Z
                           => n1711);
   U2173 : MUX2_X1 port map( A => REGISTERS_33_18_port, B => 
                           REGISTERS_34_18_port, S => n762, Z => n1712);
   U2174 : MUX2_X1 port map( A => REGISTERS_31_18_port, B => 
                           REGISTERS_32_18_port, S => n762, Z => n1713);
   U2175 : MUX2_X1 port map( A => n1713, B => n1712, S => n816, Z => n1714);
   U2176 : MUX2_X1 port map( A => REGISTERS_17_18_port, B => 
                           REGISTERS_18_18_port, S => n762, Z => n1715);
   U2177 : MUX2_X1 port map( A => REGISTERS_15_18_port, B => 
                           REGISTERS_16_18_port, S => n762, Z => n1716);
   U2178 : MUX2_X1 port map( A => n1716, B => n1715, S => n816, Z => n1717);
   U2179 : MUX2_X1 port map( A => n1717, B => n1714, S => n843, Z => n1718);
   U2180 : MUX2_X1 port map( A => n1718, B => n1711, S => n848, Z => n1719);
   U2181 : MUX2_X1 port map( A => REGISTERS_25_18_port, B => 
                           REGISTERS_26_18_port, S => n762, Z => n1720);
   U2182 : MUX2_X1 port map( A => REGISTERS_23_18_port, B => 
                           REGISTERS_24_18_port, S => n762, Z => n1721);
   U2183 : MUX2_X1 port map( A => n1721, B => n1720, S => n816, Z => n1722);
   U2184 : MUX2_X1 port map( A => REGISTERS_9_18_port, B => 
                           REGISTERS_10_18_port, S => n762, Z => n1723);
   U2185 : MUX2_X1 port map( A => REGISTERS_7_18_port, B => REGISTERS_8_18_port
                           , S => n762, Z => n1724);
   U2186 : MUX2_X1 port map( A => n1724, B => n1723, S => n816, Z => n1725);
   U2187 : MUX2_X1 port map( A => n1725, B => n1722, S => n843, Z => n1726);
   U2188 : MUX2_X1 port map( A => n1726, B => REGISTERS_39_18_port, S => n848, 
                           Z => n1727);
   U2189 : MUX2_X1 port map( A => n1727, B => n1719, S => n302, Z => n1728);
   U2190 : MUX2_X1 port map( A => n1728, B => n1709, S => n301, Z => N12223);
   U2191 : MUX2_X1 port map( A => REGISTERS_5_19_port, B => REGISTERS_6_19_port
                           , S => n761, Z => n1729);
   U2192 : MUX2_X1 port map( A => REGISTERS_3_19_port, B => REGISTERS_4_19_port
                           , S => n761, Z => n1730);
   U2193 : MUX2_X1 port map( A => n1730, B => n1729, S => n816, Z => n1731);
   U2194 : MUX2_X1 port map( A => REGISTERS_37_19_port, B => 
                           REGISTERS_38_19_port, S => n761, Z => n1732);
   U2195 : MUX2_X1 port map( A => REGISTERS_35_19_port, B => 
                           REGISTERS_36_19_port, S => n761, Z => n1733);
   U2196 : MUX2_X1 port map( A => n1733, B => n1732, S => n816, Z => n1734);
   U2197 : MUX2_X1 port map( A => REGISTERS_21_19_port, B => 
                           REGISTERS_22_19_port, S => n761, Z => n1735);
   U2198 : MUX2_X1 port map( A => REGISTERS_19_19_port, B => 
                           REGISTERS_20_19_port, S => n761, Z => n1736);
   U2199 : MUX2_X1 port map( A => n1736, B => n1735, S => n816, Z => n1737);
   U2200 : MUX2_X1 port map( A => n1737, B => n1734, S => n843, Z => n1738);
   U2201 : MUX2_X1 port map( A => n1738, B => n1731, S => n848, Z => n1739);
   U2202 : MUX2_X1 port map( A => REGISTERS_29_19_port, B => 
                           REGISTERS_30_19_port, S => n761, Z => n1740);
   U2203 : MUX2_X1 port map( A => REGISTERS_27_19_port, B => 
                           REGISTERS_28_19_port, S => n761, Z => n1741);
   U2204 : MUX2_X1 port map( A => n1741, B => n1740, S => n816, Z => n1742);
   U2205 : MUX2_X1 port map( A => REGISTERS_13_19_port, B => 
                           REGISTERS_14_19_port, S => n761, Z => n1743);
   U2206 : MUX2_X1 port map( A => REGISTERS_11_19_port, B => 
                           REGISTERS_12_19_port, S => n761, Z => n1744);
   U2207 : MUX2_X1 port map( A => n1744, B => n1743, S => n817, Z => n1745);
   U2208 : MUX2_X1 port map( A => n1745, B => n1742, S => n843, Z => n1746);
   U2209 : MUX2_X1 port map( A => n1746, B => n1739, S => n302, Z => n1747);
   U2210 : MUX2_X1 port map( A => REGISTERS_1_19_port, B => REGISTERS_2_19_port
                           , S => n761, Z => n1748);
   U2211 : MUX2_X1 port map( A => REGISTERS_0_19_port, B => n1748, S => n817, Z
                           => n1749);
   U2212 : MUX2_X1 port map( A => REGISTERS_33_19_port, B => 
                           REGISTERS_34_19_port, S => n761, Z => n1750);
   U2213 : MUX2_X1 port map( A => REGISTERS_31_19_port, B => 
                           REGISTERS_32_19_port, S => n760, Z => n1751);
   U2214 : MUX2_X1 port map( A => n1751, B => n1750, S => n817, Z => n1752);
   U2215 : MUX2_X1 port map( A => REGISTERS_17_19_port, B => 
                           REGISTERS_18_19_port, S => n760, Z => n1753);
   U2216 : MUX2_X1 port map( A => REGISTERS_15_19_port, B => 
                           REGISTERS_16_19_port, S => n760, Z => n1754);
   U2217 : MUX2_X1 port map( A => n1754, B => n1753, S => n817, Z => n1755);
   U2218 : MUX2_X1 port map( A => n1755, B => n1752, S => n843, Z => n1756);
   U2219 : MUX2_X1 port map( A => n1756, B => n1749, S => n848, Z => n1757);
   U2220 : MUX2_X1 port map( A => REGISTERS_25_19_port, B => 
                           REGISTERS_26_19_port, S => n760, Z => n1758);
   U2221 : MUX2_X1 port map( A => REGISTERS_23_19_port, B => 
                           REGISTERS_24_19_port, S => n760, Z => n1759);
   U2222 : MUX2_X1 port map( A => n1759, B => n1758, S => n817, Z => n1760);
   U2223 : MUX2_X1 port map( A => REGISTERS_9_19_port, B => 
                           REGISTERS_10_19_port, S => n760, Z => n1761);
   U2224 : MUX2_X1 port map( A => REGISTERS_7_19_port, B => REGISTERS_8_19_port
                           , S => n760, Z => n1762);
   U2225 : MUX2_X1 port map( A => n1762, B => n1761, S => n817, Z => n1763);
   U2226 : MUX2_X1 port map( A => n1763, B => n1760, S => n843, Z => n1764);
   U2227 : MUX2_X1 port map( A => n1764, B => REGISTERS_39_19_port, S => n847, 
                           Z => n1765);
   U2228 : MUX2_X1 port map( A => n1765, B => n1757, S => n302, Z => n1766);
   U2229 : MUX2_X1 port map( A => n1766, B => n1747, S => n301, Z => N12224);
   U2230 : MUX2_X1 port map( A => REGISTERS_5_20_port, B => REGISTERS_6_20_port
                           , S => n760, Z => n1767);
   U2231 : MUX2_X1 port map( A => REGISTERS_3_20_port, B => REGISTERS_4_20_port
                           , S => n760, Z => n1768);
   U2232 : MUX2_X1 port map( A => n1768, B => n1767, S => n817, Z => n1769);
   U2233 : MUX2_X1 port map( A => REGISTERS_37_20_port, B => 
                           REGISTERS_38_20_port, S => n760, Z => n1770);
   U2234 : MUX2_X1 port map( A => REGISTERS_35_20_port, B => 
                           REGISTERS_36_20_port, S => n760, Z => n1771);
   U2235 : MUX2_X1 port map( A => n1771, B => n1770, S => n817, Z => n1772);
   U2236 : MUX2_X1 port map( A => REGISTERS_21_20_port, B => 
                           REGISTERS_22_20_port, S => n759, Z => n1773);
   U2237 : MUX2_X1 port map( A => REGISTERS_19_20_port, B => 
                           REGISTERS_20_20_port, S => n759, Z => n1774);
   U2238 : MUX2_X1 port map( A => n1774, B => n1773, S => n817, Z => n1775);
   U2239 : MUX2_X1 port map( A => n1775, B => n1772, S => n843, Z => n1776);
   U2240 : MUX2_X1 port map( A => n1776, B => n1769, S => n847, Z => n1777);
   U2241 : MUX2_X1 port map( A => REGISTERS_29_20_port, B => 
                           REGISTERS_30_20_port, S => n759, Z => n1778);
   U2242 : MUX2_X1 port map( A => REGISTERS_27_20_port, B => 
                           REGISTERS_28_20_port, S => n759, Z => n1779);
   U2243 : MUX2_X1 port map( A => n1779, B => n1778, S => n817, Z => n1780);
   U2244 : MUX2_X1 port map( A => REGISTERS_13_20_port, B => 
                           REGISTERS_14_20_port, S => n759, Z => n1781);
   U2245 : MUX2_X1 port map( A => REGISTERS_11_20_port, B => 
                           REGISTERS_12_20_port, S => n759, Z => n1782);
   U2246 : MUX2_X1 port map( A => n1782, B => n1781, S => n817, Z => n1783);
   U2247 : MUX2_X1 port map( A => n1783, B => n1780, S => n843, Z => n1784);
   U2248 : MUX2_X1 port map( A => n1784, B => n1777, S => n302, Z => n1785);
   U2249 : MUX2_X1 port map( A => REGISTERS_1_20_port, B => REGISTERS_2_20_port
                           , S => n759, Z => n1786);
   U2250 : MUX2_X1 port map( A => REGISTERS_0_20_port, B => n1786, S => n817, Z
                           => n1787);
   U2251 : MUX2_X1 port map( A => REGISTERS_33_20_port, B => 
                           REGISTERS_34_20_port, S => n759, Z => n1788);
   U2252 : MUX2_X1 port map( A => REGISTERS_31_20_port, B => 
                           REGISTERS_32_20_port, S => n759, Z => n1789);
   U2253 : MUX2_X1 port map( A => n1789, B => n1788, S => n818, Z => n1790);
   U2254 : MUX2_X1 port map( A => REGISTERS_17_20_port, B => 
                           REGISTERS_18_20_port, S => n759, Z => n1791);
   U2255 : MUX2_X1 port map( A => REGISTERS_15_20_port, B => 
                           REGISTERS_16_20_port, S => n759, Z => n1792);
   U2256 : MUX2_X1 port map( A => n1792, B => n1791, S => n818, Z => n1793);
   U2257 : MUX2_X1 port map( A => n1793, B => n1790, S => n843, Z => n1794);
   U2258 : MUX2_X1 port map( A => n1794, B => n1787, S => n847, Z => n1795);
   U2259 : MUX2_X1 port map( A => REGISTERS_25_20_port, B => 
                           REGISTERS_26_20_port, S => n759, Z => n1796);
   U2260 : MUX2_X1 port map( A => REGISTERS_23_20_port, B => 
                           REGISTERS_24_20_port, S => n758, Z => n1797);
   U2261 : MUX2_X1 port map( A => n1797, B => n1796, S => n818, Z => n1798);
   U2262 : MUX2_X1 port map( A => REGISTERS_9_20_port, B => 
                           REGISTERS_10_20_port, S => n758, Z => n1799);
   U2263 : MUX2_X1 port map( A => REGISTERS_7_20_port, B => REGISTERS_8_20_port
                           , S => n758, Z => n1800);
   U2264 : MUX2_X1 port map( A => n1800, B => n1799, S => n818, Z => n1801);
   U2265 : MUX2_X1 port map( A => n1801, B => n1798, S => n843, Z => n1802);
   U2266 : MUX2_X1 port map( A => n1802, B => REGISTERS_39_20_port, S => n847, 
                           Z => n1803);
   U2267 : MUX2_X1 port map( A => n1803, B => n1795, S => n302, Z => n1804);
   U2268 : MUX2_X1 port map( A => n1804, B => n1785, S => n301, Z => N12225);
   U2269 : MUX2_X1 port map( A => REGISTERS_5_21_port, B => REGISTERS_6_21_port
                           , S => n758, Z => n1805);
   U2270 : MUX2_X1 port map( A => REGISTERS_3_21_port, B => REGISTERS_4_21_port
                           , S => n758, Z => n1806);
   U2271 : MUX2_X1 port map( A => n1806, B => n1805, S => n818, Z => n1807);
   U2272 : MUX2_X1 port map( A => REGISTERS_37_21_port, B => 
                           REGISTERS_38_21_port, S => n758, Z => n1808);
   U2273 : MUX2_X1 port map( A => REGISTERS_35_21_port, B => 
                           REGISTERS_36_21_port, S => n758, Z => n1809);
   U2274 : MUX2_X1 port map( A => n1809, B => n1808, S => n818, Z => n1810);
   U2275 : MUX2_X1 port map( A => REGISTERS_21_21_port, B => 
                           REGISTERS_22_21_port, S => n758, Z => n1811);
   U2276 : MUX2_X1 port map( A => REGISTERS_19_21_port, B => 
                           REGISTERS_20_21_port, S => n758, Z => n1812);
   U2277 : MUX2_X1 port map( A => n1812, B => n1811, S => n818, Z => n1813);
   U2278 : MUX2_X1 port map( A => n1813, B => n1810, S => n843, Z => n1814);
   U2279 : MUX2_X1 port map( A => n1814, B => n1807, S => n847, Z => n1815);
   U2280 : MUX2_X1 port map( A => REGISTERS_29_21_port, B => 
                           REGISTERS_30_21_port, S => n758, Z => n1816);
   U2281 : MUX2_X1 port map( A => REGISTERS_27_21_port, B => 
                           REGISTERS_28_21_port, S => n758, Z => n1817);
   U2282 : MUX2_X1 port map( A => n1817, B => n1816, S => n818, Z => n1818);
   U2283 : MUX2_X1 port map( A => REGISTERS_13_21_port, B => 
                           REGISTERS_14_21_port, S => n758, Z => n1819);
   U2284 : MUX2_X1 port map( A => REGISTERS_11_21_port, B => 
                           REGISTERS_12_21_port, S => n757, Z => n1820);
   U2285 : MUX2_X1 port map( A => n1820, B => n1819, S => n818, Z => n1821);
   U2286 : MUX2_X1 port map( A => n1821, B => n1818, S => n843, Z => n1822);
   U2287 : MUX2_X1 port map( A => n1822, B => n1815, S => n302, Z => n1823);
   U2288 : MUX2_X1 port map( A => REGISTERS_1_21_port, B => REGISTERS_2_21_port
                           , S => n757, Z => n1824);
   U2289 : MUX2_X1 port map( A => REGISTERS_0_21_port, B => n1824, S => n818, Z
                           => n1825);
   U2290 : MUX2_X1 port map( A => REGISTERS_33_21_port, B => 
                           REGISTERS_34_21_port, S => n757, Z => n1826);
   U2291 : MUX2_X1 port map( A => REGISTERS_31_21_port, B => 
                           REGISTERS_32_21_port, S => n757, Z => n1827);
   U2292 : MUX2_X1 port map( A => n1827, B => n1826, S => n818, Z => n1828);
   U2293 : MUX2_X1 port map( A => REGISTERS_17_21_port, B => 
                           REGISTERS_18_21_port, S => n757, Z => n1829);
   U2294 : MUX2_X1 port map( A => REGISTERS_15_21_port, B => 
                           REGISTERS_16_21_port, S => n757, Z => n1830);
   U2295 : MUX2_X1 port map( A => n1830, B => n1829, S => n818, Z => n1831);
   U2296 : MUX2_X1 port map( A => n1831, B => n1828, S => n843, Z => n1832);
   U2297 : MUX2_X1 port map( A => n1832, B => n1825, S => n847, Z => n1833);
   U2298 : MUX2_X1 port map( A => REGISTERS_25_21_port, B => 
                           REGISTERS_26_21_port, S => n757, Z => n1834);
   U2299 : MUX2_X1 port map( A => REGISTERS_23_21_port, B => 
                           REGISTERS_24_21_port, S => n757, Z => n1835);
   U2300 : MUX2_X1 port map( A => n1835, B => n1834, S => n819, Z => n1836);
   U2301 : MUX2_X1 port map( A => REGISTERS_9_21_port, B => 
                           REGISTERS_10_21_port, S => n757, Z => n1837);
   U2302 : MUX2_X1 port map( A => REGISTERS_7_21_port, B => REGISTERS_8_21_port
                           , S => n757, Z => n1838);
   U2303 : MUX2_X1 port map( A => n1838, B => n1837, S => n819, Z => n1839);
   U2304 : MUX2_X1 port map( A => n1839, B => n1836, S => n843, Z => n1840);
   U2305 : MUX2_X1 port map( A => n1840, B => REGISTERS_39_21_port, S => n847, 
                           Z => n1841);
   U2306 : MUX2_X1 port map( A => n1841, B => n1833, S => n302, Z => n1842);
   U2307 : MUX2_X1 port map( A => n1842, B => n1823, S => n301, Z => N12226);
   U2308 : MUX2_X1 port map( A => REGISTERS_5_22_port, B => REGISTERS_6_22_port
                           , S => n757, Z => n1843);
   U2309 : MUX2_X1 port map( A => REGISTERS_3_22_port, B => REGISTERS_4_22_port
                           , S => n757, Z => n1844);
   U2310 : MUX2_X1 port map( A => n1844, B => n1843, S => n819, Z => n1845);
   U2311 : MUX2_X1 port map( A => REGISTERS_37_22_port, B => 
                           REGISTERS_38_22_port, S => n756, Z => n1846);
   U2312 : MUX2_X1 port map( A => REGISTERS_35_22_port, B => 
                           REGISTERS_36_22_port, S => n756, Z => n1847);
   U2313 : MUX2_X1 port map( A => n1847, B => n1846, S => n819, Z => n1848);
   U2314 : MUX2_X1 port map( A => REGISTERS_21_22_port, B => 
                           REGISTERS_22_22_port, S => n756, Z => n1849);
   U2315 : MUX2_X1 port map( A => REGISTERS_19_22_port, B => 
                           REGISTERS_20_22_port, S => n756, Z => n1850);
   U2316 : MUX2_X1 port map( A => n1850, B => n1849, S => n819, Z => n1851);
   U2317 : MUX2_X1 port map( A => n1851, B => n1848, S => n843, Z => n1852);
   U2318 : MUX2_X1 port map( A => n1852, B => n1845, S => n847, Z => n1853);
   U2319 : MUX2_X1 port map( A => REGISTERS_29_22_port, B => 
                           REGISTERS_30_22_port, S => n756, Z => n1854);
   U2320 : MUX2_X1 port map( A => REGISTERS_27_22_port, B => 
                           REGISTERS_28_22_port, S => n756, Z => n1855);
   U2321 : MUX2_X1 port map( A => n1855, B => n1854, S => n819, Z => n1856);
   U2322 : MUX2_X1 port map( A => REGISTERS_13_22_port, B => 
                           REGISTERS_14_22_port, S => n756, Z => n1857);
   U2323 : MUX2_X1 port map( A => REGISTERS_11_22_port, B => 
                           REGISTERS_12_22_port, S => n756, Z => n1858);
   U2324 : MUX2_X1 port map( A => n1858, B => n1857, S => n819, Z => n1859);
   U2325 : MUX2_X1 port map( A => n1859, B => n1856, S => n843, Z => n1860);
   U2326 : MUX2_X1 port map( A => n1860, B => n1853, S => n302, Z => n1861);
   U2327 : MUX2_X1 port map( A => REGISTERS_1_22_port, B => REGISTERS_2_22_port
                           , S => n756, Z => n1862);
   U2328 : MUX2_X1 port map( A => REGISTERS_0_22_port, B => n1862, S => n819, Z
                           => n1863);
   U2329 : MUX2_X1 port map( A => REGISTERS_33_22_port, B => 
                           REGISTERS_34_22_port, S => n756, Z => n1864);
   U2330 : MUX2_X1 port map( A => REGISTERS_31_22_port, B => 
                           REGISTERS_32_22_port, S => n756, Z => n1865);
   U2331 : MUX2_X1 port map( A => n1865, B => n1864, S => n819, Z => n1866);
   U2332 : MUX2_X1 port map( A => REGISTERS_17_22_port, B => 
                           REGISTERS_18_22_port, S => n756, Z => n1867);
   U2333 : MUX2_X1 port map( A => REGISTERS_15_22_port, B => 
                           REGISTERS_16_22_port, S => n755, Z => n1868);
   U2334 : MUX2_X1 port map( A => n1868, B => n1867, S => n819, Z => n1869);
   U2335 : MUX2_X1 port map( A => n1869, B => n1866, S => n842, Z => n1870);
   U2336 : MUX2_X1 port map( A => n1870, B => n1863, S => n847, Z => n1871);
   U2337 : MUX2_X1 port map( A => REGISTERS_25_22_port, B => 
                           REGISTERS_26_22_port, S => n755, Z => n1872);
   U2338 : MUX2_X1 port map( A => REGISTERS_23_22_port, B => 
                           REGISTERS_24_22_port, S => n755, Z => n1873);
   U2339 : MUX2_X1 port map( A => n1873, B => n1872, S => n819, Z => n1874);
   U2340 : MUX2_X1 port map( A => REGISTERS_9_22_port, B => 
                           REGISTERS_10_22_port, S => n755, Z => n1875);
   U2341 : MUX2_X1 port map( A => REGISTERS_7_22_port, B => REGISTERS_8_22_port
                           , S => n755, Z => n1876);
   U2342 : MUX2_X1 port map( A => n1876, B => n1875, S => n819, Z => n1877);
   U2343 : MUX2_X1 port map( A => n1877, B => n1874, S => n842, Z => n1878);
   U2344 : MUX2_X1 port map( A => n1878, B => REGISTERS_39_22_port, S => n847, 
                           Z => n1879);
   U2345 : MUX2_X1 port map( A => n1879, B => n1871, S => n302, Z => n1880);
   U2346 : MUX2_X1 port map( A => n1880, B => n1861, S => n301, Z => N12227);
   U2347 : MUX2_X1 port map( A => REGISTERS_5_23_port, B => REGISTERS_6_23_port
                           , S => n755, Z => n1881);
   U2348 : MUX2_X1 port map( A => REGISTERS_3_23_port, B => REGISTERS_4_23_port
                           , S => n755, Z => n1882);
   U2349 : MUX2_X1 port map( A => n1882, B => n1881, S => n820, Z => n1883);
   U2350 : MUX2_X1 port map( A => REGISTERS_37_23_port, B => 
                           REGISTERS_38_23_port, S => n755, Z => n1884);
   U2351 : MUX2_X1 port map( A => REGISTERS_35_23_port, B => 
                           REGISTERS_36_23_port, S => n755, Z => n1885);
   U2352 : MUX2_X1 port map( A => n1885, B => n1884, S => n820, Z => n1886);
   U2353 : MUX2_X1 port map( A => REGISTERS_21_23_port, B => 
                           REGISTERS_22_23_port, S => n755, Z => n1887);
   U2354 : MUX2_X1 port map( A => REGISTERS_19_23_port, B => 
                           REGISTERS_20_23_port, S => n755, Z => n1888);
   U2355 : MUX2_X1 port map( A => n1888, B => n1887, S => n820, Z => n1889);
   U2356 : MUX2_X1 port map( A => n1889, B => n1886, S => n842, Z => n1890);
   U2357 : MUX2_X1 port map( A => n1890, B => n1883, S => n847, Z => n1891);
   U2358 : MUX2_X1 port map( A => REGISTERS_29_23_port, B => 
                           REGISTERS_30_23_port, S => n755, Z => n1892);
   U2359 : MUX2_X1 port map( A => REGISTERS_27_23_port, B => 
                           REGISTERS_28_23_port, S => n754, Z => n1893);
   U2360 : MUX2_X1 port map( A => n1893, B => n1892, S => n820, Z => n1894);
   U2361 : MUX2_X1 port map( A => REGISTERS_13_23_port, B => 
                           REGISTERS_14_23_port, S => n754, Z => n1895);
   U2362 : MUX2_X1 port map( A => REGISTERS_11_23_port, B => 
                           REGISTERS_12_23_port, S => n754, Z => n1896);
   U2363 : MUX2_X1 port map( A => n1896, B => n1895, S => n820, Z => n1897);
   U2364 : MUX2_X1 port map( A => n1897, B => n1894, S => n842, Z => n1898);
   U2365 : MUX2_X1 port map( A => n1898, B => n1891, S => n302, Z => n1899);
   U2366 : MUX2_X1 port map( A => REGISTERS_1_23_port, B => REGISTERS_2_23_port
                           , S => n754, Z => n1900);
   U2367 : MUX2_X1 port map( A => REGISTERS_0_23_port, B => n1900, S => n820, Z
                           => n1901);
   U2368 : MUX2_X1 port map( A => REGISTERS_33_23_port, B => 
                           REGISTERS_34_23_port, S => n754, Z => n1902);
   U2369 : MUX2_X1 port map( A => REGISTERS_31_23_port, B => 
                           REGISTERS_32_23_port, S => n754, Z => n1903);
   U2370 : MUX2_X1 port map( A => n1903, B => n1902, S => n820, Z => n1904);
   U2371 : MUX2_X1 port map( A => REGISTERS_17_23_port, B => 
                           REGISTERS_18_23_port, S => n754, Z => n1905);
   U2372 : MUX2_X1 port map( A => REGISTERS_15_23_port, B => 
                           REGISTERS_16_23_port, S => n754, Z => n1906);
   U2373 : MUX2_X1 port map( A => n1906, B => n1905, S => n820, Z => n1907);
   U2374 : MUX2_X1 port map( A => n1907, B => n1904, S => n842, Z => n1908);
   U2375 : MUX2_X1 port map( A => n1908, B => n1901, S => n847, Z => n1909);
   U2376 : MUX2_X1 port map( A => REGISTERS_25_23_port, B => 
                           REGISTERS_26_23_port, S => n754, Z => n1910);
   U2377 : MUX2_X1 port map( A => REGISTERS_23_23_port, B => 
                           REGISTERS_24_23_port, S => n754, Z => n1911);
   U2378 : MUX2_X1 port map( A => n1911, B => n1910, S => n820, Z => n1912);
   U2379 : MUX2_X1 port map( A => REGISTERS_9_23_port, B => 
                           REGISTERS_10_23_port, S => n760, Z => n1913);
   U2380 : MUX2_X1 port map( A => REGISTERS_7_23_port, B => REGISTERS_8_23_port
                           , S => n779, Z => n1914);
   U2381 : MUX2_X1 port map( A => n1914, B => n1913, S => n820, Z => n1915);
   U2382 : MUX2_X1 port map( A => n1915, B => n1912, S => n842, Z => n1916);
   U2383 : MUX2_X1 port map( A => n1916, B => REGISTERS_39_23_port, S => n847, 
                           Z => n1917);
   U2384 : MUX2_X1 port map( A => n1917, B => n1909, S => n302, Z => n1918);
   U2385 : MUX2_X1 port map( A => n1918, B => n1899, S => n301, Z => N12228);
   U2386 : MUX2_X1 port map( A => REGISTERS_5_24_port, B => REGISTERS_6_24_port
                           , S => n779, Z => n1919);
   U2387 : MUX2_X1 port map( A => REGISTERS_3_24_port, B => REGISTERS_4_24_port
                           , S => n779, Z => n1920);
   U2388 : MUX2_X1 port map( A => n1920, B => n1919, S => n820, Z => n1921);
   U2389 : MUX2_X1 port map( A => REGISTERS_37_24_port, B => 
                           REGISTERS_38_24_port, S => n779, Z => n1922);
   U2390 : MUX2_X1 port map( A => REGISTERS_35_24_port, B => 
                           REGISTERS_36_24_port, S => n779, Z => n1923);
   U2391 : MUX2_X1 port map( A => n1923, B => n1922, S => n821, Z => n1924);
   U2392 : MUX2_X1 port map( A => REGISTERS_21_24_port, B => 
                           REGISTERS_22_24_port, S => n778, Z => n1925);
   U2393 : MUX2_X1 port map( A => REGISTERS_19_24_port, B => 
                           REGISTERS_20_24_port, S => n778, Z => n1926);
   U2394 : MUX2_X1 port map( A => n1926, B => n1925, S => n821, Z => n1927);
   U2395 : MUX2_X1 port map( A => n1927, B => n1924, S => n842, Z => n1928);
   U2396 : MUX2_X1 port map( A => n1928, B => n1921, S => n847, Z => n1929);
   U2397 : MUX2_X1 port map( A => REGISTERS_29_24_port, B => 
                           REGISTERS_30_24_port, S => n778, Z => n1930);
   U2398 : MUX2_X1 port map( A => REGISTERS_27_24_port, B => 
                           REGISTERS_28_24_port, S => n778, Z => n1931);
   U2399 : MUX2_X1 port map( A => n1931, B => n1930, S => n821, Z => n1932);
   U2400 : MUX2_X1 port map( A => REGISTERS_13_24_port, B => 
                           REGISTERS_14_24_port, S => n778, Z => n1933);
   U2401 : MUX2_X1 port map( A => REGISTERS_11_24_port, B => 
                           REGISTERS_12_24_port, S => n778, Z => n1934);
   U2402 : MUX2_X1 port map( A => n1934, B => n1933, S => n821, Z => n1935);
   U2403 : MUX2_X1 port map( A => n1935, B => n1932, S => n842, Z => n1936);
   U2404 : MUX2_X1 port map( A => n1936, B => n1929, S => n302, Z => n1937);
   U2405 : MUX2_X1 port map( A => REGISTERS_1_24_port, B => REGISTERS_2_24_port
                           , S => n778, Z => n1938);
   U2406 : MUX2_X1 port map( A => REGISTERS_0_24_port, B => n1938, S => n821, Z
                           => n1939);
   U2407 : MUX2_X1 port map( A => REGISTERS_33_24_port, B => 
                           REGISTERS_34_24_port, S => n778, Z => n1940);
   U2408 : MUX2_X1 port map( A => REGISTERS_31_24_port, B => 
                           REGISTERS_32_24_port, S => n778, Z => n1941);
   U2409 : MUX2_X1 port map( A => n1941, B => n1940, S => n821, Z => n1942);
   U2410 : MUX2_X1 port map( A => REGISTERS_17_24_port, B => 
                           REGISTERS_18_24_port, S => n778, Z => n1943);
   U2411 : MUX2_X1 port map( A => REGISTERS_15_24_port, B => 
                           REGISTERS_16_24_port, S => n778, Z => n1944);
   U2412 : MUX2_X1 port map( A => n1944, B => n1943, S => n821, Z => n1945);
   U2413 : MUX2_X1 port map( A => n1945, B => n1942, S => n842, Z => n1946);
   U2414 : MUX2_X1 port map( A => n1946, B => n1939, S => n847, Z => n1947);
   U2415 : MUX2_X1 port map( A => REGISTERS_25_24_port, B => 
                           REGISTERS_26_24_port, S => n778, Z => n1948);
   U2416 : MUX2_X1 port map( A => REGISTERS_23_24_port, B => 
                           REGISTERS_24_24_port, S => n777, Z => n1949);
   U2417 : MUX2_X1 port map( A => n1949, B => n1948, S => n821, Z => n1950);
   U2418 : MUX2_X1 port map( A => REGISTERS_9_24_port, B => 
                           REGISTERS_10_24_port, S => n777, Z => n1951);
   U2419 : MUX2_X1 port map( A => REGISTERS_7_24_port, B => REGISTERS_8_24_port
                           , S => n777, Z => n1952);
   U2420 : MUX2_X1 port map( A => n1952, B => n1951, S => n821, Z => n1953);
   U2421 : MUX2_X1 port map( A => n1953, B => n1950, S => n842, Z => n1954);
   U2422 : MUX2_X1 port map( A => n1954, B => REGISTERS_39_24_port, S => n847, 
                           Z => n1955);
   U2423 : MUX2_X1 port map( A => n1955, B => n1947, S => n302, Z => n1956);
   U2424 : MUX2_X1 port map( A => n1956, B => n1937, S => n301, Z => N12229);
   U2425 : MUX2_X1 port map( A => REGISTERS_5_25_port, B => REGISTERS_6_25_port
                           , S => n777, Z => n1957);
   U2426 : MUX2_X1 port map( A => REGISTERS_3_25_port, B => REGISTERS_4_25_port
                           , S => n777, Z => n1958);
   U2427 : MUX2_X1 port map( A => n1958, B => n1957, S => n821, Z => n1959);
   U2428 : MUX2_X1 port map( A => REGISTERS_37_25_port, B => 
                           REGISTERS_38_25_port, S => n777, Z => n1960);
   U2429 : MUX2_X1 port map( A => REGISTERS_35_25_port, B => 
                           REGISTERS_36_25_port, S => n777, Z => n1961);
   U2430 : MUX2_X1 port map( A => n1961, B => n1960, S => n821, Z => n1962);
   U2431 : MUX2_X1 port map( A => REGISTERS_21_25_port, B => 
                           REGISTERS_22_25_port, S => n777, Z => n1963);
   U2432 : MUX2_X1 port map( A => REGISTERS_19_25_port, B => 
                           REGISTERS_20_25_port, S => n777, Z => n1964);
   U2433 : MUX2_X1 port map( A => n1964, B => n1963, S => n821, Z => n1965);
   U2434 : MUX2_X1 port map( A => n1965, B => n1962, S => n842, Z => n1966);
   U2435 : MUX2_X1 port map( A => n1966, B => n1959, S => n847, Z => n1967);
   U2436 : MUX2_X1 port map( A => REGISTERS_29_25_port, B => 
                           REGISTERS_30_25_port, S => n777, Z => n1968);
   U2437 : MUX2_X1 port map( A => REGISTERS_27_25_port, B => 
                           REGISTERS_28_25_port, S => n777, Z => n1969);
   U2438 : MUX2_X1 port map( A => n1969, B => n1968, S => n822, Z => n1970);
   U2439 : MUX2_X1 port map( A => REGISTERS_13_25_port, B => 
                           REGISTERS_14_25_port, S => n777, Z => n1971);
   U2440 : MUX2_X1 port map( A => REGISTERS_11_25_port, B => 
                           REGISTERS_12_25_port, S => n776, Z => n1972);
   U2441 : MUX2_X1 port map( A => n1972, B => n1971, S => n822, Z => n1973);
   U2442 : MUX2_X1 port map( A => n1973, B => n1970, S => n842, Z => n1974);
   U2443 : MUX2_X1 port map( A => n1974, B => n1967, S => n302, Z => n1975);
   U2444 : MUX2_X1 port map( A => REGISTERS_1_25_port, B => REGISTERS_2_25_port
                           , S => n776, Z => n1976);
   U2445 : MUX2_X1 port map( A => REGISTERS_0_25_port, B => n1976, S => n822, Z
                           => n1977);
   U2446 : MUX2_X1 port map( A => REGISTERS_33_25_port, B => 
                           REGISTERS_34_25_port, S => n776, Z => n1978);
   U2447 : MUX2_X1 port map( A => REGISTERS_31_25_port, B => 
                           REGISTERS_32_25_port, S => n776, Z => n1979);
   U2448 : MUX2_X1 port map( A => n1979, B => n1978, S => n822, Z => n1980);
   U2449 : MUX2_X1 port map( A => REGISTERS_17_25_port, B => 
                           REGISTERS_18_25_port, S => n776, Z => n1981);
   U2450 : MUX2_X1 port map( A => REGISTERS_15_25_port, B => 
                           REGISTERS_16_25_port, S => n776, Z => n1982);
   U2451 : MUX2_X1 port map( A => n1982, B => n1981, S => n822, Z => n1983);
   U2452 : MUX2_X1 port map( A => n1983, B => n1980, S => n842, Z => n1984);
   U2453 : MUX2_X1 port map( A => n1984, B => n1977, S => n847, Z => n1985);
   U2454 : MUX2_X1 port map( A => REGISTERS_25_25_port, B => 
                           REGISTERS_26_25_port, S => n776, Z => n1986);
   U2455 : MUX2_X1 port map( A => REGISTERS_23_25_port, B => 
                           REGISTERS_24_25_port, S => n776, Z => n1987);
   U2456 : MUX2_X1 port map( A => n1987, B => n1986, S => n822, Z => n1988);
   U2457 : MUX2_X1 port map( A => REGISTERS_9_25_port, B => 
                           REGISTERS_10_25_port, S => n776, Z => n1989);
   U2458 : MUX2_X1 port map( A => REGISTERS_7_25_port, B => REGISTERS_8_25_port
                           , S => n776, Z => n1990);
   U2459 : MUX2_X1 port map( A => n1990, B => n1989, S => n822, Z => n1991);
   U2460 : MUX2_X1 port map( A => n1991, B => n1988, S => n842, Z => n1992);
   U2461 : MUX2_X1 port map( A => n1992, B => REGISTERS_39_25_port, S => n847, 
                           Z => n1993);
   U2462 : MUX2_X1 port map( A => n1993, B => n1985, S => n302, Z => n1994);
   U2463 : MUX2_X1 port map( A => n1994, B => n1975, S => n301, Z => N12230);
   U2464 : MUX2_X1 port map( A => REGISTERS_5_26_port, B => REGISTERS_6_26_port
                           , S => n776, Z => n1995);
   U2465 : MUX2_X1 port map( A => REGISTERS_3_26_port, B => REGISTERS_4_26_port
                           , S => n776, Z => n1996);
   U2466 : MUX2_X1 port map( A => n1996, B => n1995, S => n822, Z => n1997);
   U2467 : MUX2_X1 port map( A => REGISTERS_37_26_port, B => 
                           REGISTERS_38_26_port, S => n775, Z => n1998);
   U2468 : MUX2_X1 port map( A => REGISTERS_35_26_port, B => 
                           REGISTERS_36_26_port, S => n775, Z => n1999);
   U2469 : MUX2_X1 port map( A => n1999, B => n1998, S => n822, Z => n2000);
   U2470 : MUX2_X1 port map( A => REGISTERS_21_26_port, B => 
                           REGISTERS_22_26_port, S => n775, Z => n2001);
   U2471 : MUX2_X1 port map( A => REGISTERS_19_26_port, B => 
                           REGISTERS_20_26_port, S => n775, Z => n2002);
   U2472 : MUX2_X1 port map( A => n2002, B => n2001, S => n822, Z => n2003);
   U2473 : MUX2_X1 port map( A => n2003, B => n2000, S => n842, Z => n2004);
   U2474 : MUX2_X1 port map( A => n2004, B => n1997, S => n847, Z => n2005);
   U2475 : MUX2_X1 port map( A => REGISTERS_29_26_port, B => 
                           REGISTERS_30_26_port, S => n775, Z => n2006);
   U2476 : MUX2_X1 port map( A => REGISTERS_27_26_port, B => 
                           REGISTERS_28_26_port, S => n775, Z => n2007);
   U2477 : MUX2_X1 port map( A => n2007, B => n2006, S => n822, Z => n2008);
   U2478 : MUX2_X1 port map( A => REGISTERS_13_26_port, B => 
                           REGISTERS_14_26_port, S => n775, Z => n2009);
   U2479 : MUX2_X1 port map( A => REGISTERS_11_26_port, B => 
                           REGISTERS_12_26_port, S => n775, Z => n2010);
   U2480 : MUX2_X1 port map( A => n2010, B => n2009, S => n822, Z => n2011);
   U2481 : MUX2_X1 port map( A => n2011, B => n2008, S => n842, Z => n2012);
   U2482 : MUX2_X1 port map( A => n2012, B => n2005, S => n302, Z => n2013);
   U2483 : MUX2_X1 port map( A => REGISTERS_1_26_port, B => REGISTERS_2_26_port
                           , S => n775, Z => n2014);
   U2484 : MUX2_X1 port map( A => REGISTERS_0_26_port, B => n2014, S => n823, Z
                           => n2015);
   U2485 : MUX2_X1 port map( A => REGISTERS_33_26_port, B => 
                           REGISTERS_34_26_port, S => n775, Z => n2016);
   U2486 : MUX2_X1 port map( A => REGISTERS_31_26_port, B => 
                           REGISTERS_32_26_port, S => n775, Z => n2017);
   U2487 : MUX2_X1 port map( A => n2017, B => n2016, S => n823, Z => n2018);
   U2488 : MUX2_X1 port map( A => REGISTERS_17_26_port, B => 
                           REGISTERS_18_26_port, S => n775, Z => n2019);
   U2489 : MUX2_X1 port map( A => REGISTERS_15_26_port, B => 
                           REGISTERS_16_26_port, S => n774, Z => n2020);
   U2490 : MUX2_X1 port map( A => n2020, B => n2019, S => n823, Z => n2021);
   U2491 : MUX2_X1 port map( A => n2021, B => n2018, S => n842, Z => n2022);
   U2492 : MUX2_X1 port map( A => n2022, B => n2015, S => n847, Z => n2023);
   U2493 : MUX2_X1 port map( A => REGISTERS_25_26_port, B => 
                           REGISTERS_26_26_port, S => n774, Z => n2024);
   U2494 : MUX2_X1 port map( A => REGISTERS_23_26_port, B => 
                           REGISTERS_24_26_port, S => n774, Z => n2025);
   U2495 : MUX2_X1 port map( A => n2025, B => n2024, S => n823, Z => n2026);
   U2496 : MUX2_X1 port map( A => REGISTERS_9_26_port, B => 
                           REGISTERS_10_26_port, S => n774, Z => n2027);
   U2497 : MUX2_X1 port map( A => REGISTERS_7_26_port, B => REGISTERS_8_26_port
                           , S => n774, Z => n2028);
   U2498 : MUX2_X1 port map( A => n2028, B => n2027, S => n823, Z => n2029);
   U2499 : MUX2_X1 port map( A => n2029, B => n2026, S => n842, Z => n2030);
   U2500 : MUX2_X1 port map( A => n2030, B => REGISTERS_39_26_port, S => n847, 
                           Z => n2031);
   U2501 : MUX2_X1 port map( A => n2031, B => n2023, S => n302, Z => n2032);
   U2502 : MUX2_X1 port map( A => n2032, B => n2013, S => n301, Z => N12231);
   U2503 : MUX2_X1 port map( A => REGISTERS_5_27_port, B => REGISTERS_6_27_port
                           , S => n774, Z => n2033);
   U2504 : MUX2_X1 port map( A => REGISTERS_3_27_port, B => REGISTERS_4_27_port
                           , S => n774, Z => n2034);
   U2505 : MUX2_X1 port map( A => n2034, B => n2033, S => n823, Z => n2035);
   U2506 : MUX2_X1 port map( A => REGISTERS_37_27_port, B => 
                           REGISTERS_38_27_port, S => n774, Z => n2036);
   U2507 : MUX2_X1 port map( A => REGISTERS_35_27_port, B => 
                           REGISTERS_36_27_port, S => n774, Z => n2037);
   U2508 : MUX2_X1 port map( A => n2037, B => n2036, S => n823, Z => n2038);
   U2509 : MUX2_X1 port map( A => REGISTERS_21_27_port, B => 
                           REGISTERS_22_27_port, S => n774, Z => n2039);
   U2510 : MUX2_X1 port map( A => REGISTERS_19_27_port, B => 
                           REGISTERS_20_27_port, S => n774, Z => n2040);
   U2511 : MUX2_X1 port map( A => n2040, B => n2039, S => n823, Z => n2041);
   U2512 : MUX2_X1 port map( A => n2041, B => n2038, S => n842, Z => n2042);
   U2513 : MUX2_X1 port map( A => n2042, B => n2035, S => n847, Z => n2043);
   U2514 : MUX2_X1 port map( A => REGISTERS_29_27_port, B => 
                           REGISTERS_30_27_port, S => n774, Z => n2044);
   U2515 : MUX2_X1 port map( A => REGISTERS_27_27_port, B => 
                           REGISTERS_28_27_port, S => n773, Z => n2045);
   U2516 : MUX2_X1 port map( A => n2045, B => n2044, S => n823, Z => n2046);
   U2517 : MUX2_X1 port map( A => REGISTERS_13_27_port, B => 
                           REGISTERS_14_27_port, S => n773, Z => n2047);
   U2518 : MUX2_X1 port map( A => REGISTERS_11_27_port, B => 
                           REGISTERS_12_27_port, S => n773, Z => n2048);
   U2519 : MUX2_X1 port map( A => n2048, B => n2047, S => n823, Z => n2049);
   U2520 : MUX2_X1 port map( A => n2049, B => n2046, S => n842, Z => n2050);
   U2521 : MUX2_X1 port map( A => n2050, B => n2043, S => n302, Z => n2051);
   U2522 : MUX2_X1 port map( A => REGISTERS_1_27_port, B => REGISTERS_2_27_port
                           , S => n773, Z => n2052);
   U2523 : MUX2_X1 port map( A => REGISTERS_0_27_port, B => n2052, S => n823, Z
                           => n2053);
   U2524 : MUX2_X1 port map( A => REGISTERS_33_27_port, B => 
                           REGISTERS_34_27_port, S => n773, Z => n2054);
   U2525 : MUX2_X1 port map( A => REGISTERS_31_27_port, B => 
                           REGISTERS_32_27_port, S => n773, Z => n2055);
   U2526 : MUX2_X1 port map( A => n2055, B => n2054, S => n823, Z => n2056);
   U2527 : MUX2_X1 port map( A => REGISTERS_17_27_port, B => 
                           REGISTERS_18_27_port, S => n773, Z => n2057);
   U2528 : MUX2_X1 port map( A => REGISTERS_15_27_port, B => 
                           REGISTERS_16_27_port, S => n773, Z => n2058);
   U2529 : MUX2_X1 port map( A => n2058, B => n2057, S => n824, Z => n2059);
   U2530 : MUX2_X1 port map( A => n2059, B => n2056, S => n842, Z => n2060);
   U2531 : MUX2_X1 port map( A => n2060, B => n2053, S => n847, Z => n2061);
   U2532 : MUX2_X1 port map( A => REGISTERS_25_27_port, B => 
                           REGISTERS_26_27_port, S => n773, Z => n2062);
   U2533 : MUX2_X1 port map( A => REGISTERS_23_27_port, B => 
                           REGISTERS_24_27_port, S => n773, Z => n2063);
   U2534 : MUX2_X1 port map( A => n2063, B => n2062, S => n824, Z => n2064);
   U2535 : MUX2_X1 port map( A => REGISTERS_9_27_port, B => 
                           REGISTERS_10_27_port, S => n773, Z => n2065);
   U2536 : MUX2_X1 port map( A => REGISTERS_7_27_port, B => REGISTERS_8_27_port
                           , S => n772, Z => n2066);
   U2537 : MUX2_X1 port map( A => n2066, B => n2065, S => n824, Z => n2067);
   U2538 : MUX2_X1 port map( A => n2067, B => n2064, S => n842, Z => n2068);
   U2539 : MUX2_X1 port map( A => n2068, B => REGISTERS_39_27_port, S => n847, 
                           Z => n2069);
   U2540 : MUX2_X1 port map( A => n2069, B => n2061, S => n302, Z => n2070);
   U2541 : MUX2_X1 port map( A => n2070, B => n2051, S => n301, Z => N12232);
   U2542 : MUX2_X1 port map( A => REGISTERS_5_28_port, B => REGISTERS_6_28_port
                           , S => n772, Z => n2071);
   U2543 : MUX2_X1 port map( A => REGISTERS_3_28_port, B => REGISTERS_4_28_port
                           , S => n772, Z => n2072);
   U2544 : MUX2_X1 port map( A => n2072, B => n2071, S => n824, Z => n2073);
   U2545 : MUX2_X1 port map( A => REGISTERS_37_28_port, B => 
                           REGISTERS_38_28_port, S => n772, Z => n2074);
   U2546 : MUX2_X1 port map( A => REGISTERS_35_28_port, B => 
                           REGISTERS_36_28_port, S => n772, Z => n2075);
   U2547 : MUX2_X1 port map( A => n2075, B => n2074, S => n824, Z => n2076);
   U2548 : MUX2_X1 port map( A => REGISTERS_21_28_port, B => 
                           REGISTERS_22_28_port, S => n772, Z => n2077);
   U2549 : MUX2_X1 port map( A => REGISTERS_19_28_port, B => 
                           REGISTERS_20_28_port, S => n772, Z => n2078);
   U2550 : MUX2_X1 port map( A => n2078, B => n2077, S => n824, Z => n2079);
   U2551 : MUX2_X1 port map( A => n2079, B => n2076, S => n842, Z => n2080);
   U2552 : MUX2_X1 port map( A => n2080, B => n2073, S => n847, Z => n2081);
   U2553 : MUX2_X1 port map( A => REGISTERS_29_28_port, B => 
                           REGISTERS_30_28_port, S => n772, Z => n2082);
   U2554 : MUX2_X1 port map( A => REGISTERS_27_28_port, B => 
                           REGISTERS_28_28_port, S => n772, Z => n2083);
   U2555 : MUX2_X1 port map( A => n2083, B => n2082, S => n824, Z => n2084);
   U2556 : MUX2_X1 port map( A => REGISTERS_13_28_port, B => 
                           REGISTERS_14_28_port, S => n772, Z => n2085);
   U2557 : MUX2_X1 port map( A => REGISTERS_11_28_port, B => 
                           REGISTERS_12_28_port, S => n772, Z => n2086);
   U2558 : MUX2_X1 port map( A => n2086, B => n2085, S => n824, Z => n2087);
   U2559 : MUX2_X1 port map( A => n2087, B => n2084, S => n842, Z => n2088);
   U2560 : MUX2_X1 port map( A => n2088, B => n2081, S => n302, Z => n2089);
   U2561 : MUX2_X1 port map( A => REGISTERS_1_28_port, B => REGISTERS_2_28_port
                           , S => n772, Z => n2090);
   U2562 : MUX2_X1 port map( A => REGISTERS_0_28_port, B => n2090, S => n824, Z
                           => n2091);
   U2563 : MUX2_X1 port map( A => REGISTERS_33_28_port, B => 
                           REGISTERS_34_28_port, S => n771, Z => n2092);
   U2564 : MUX2_X1 port map( A => REGISTERS_31_28_port, B => 
                           REGISTERS_32_28_port, S => n771, Z => n2093);
   U2565 : MUX2_X1 port map( A => n2093, B => n2092, S => n824, Z => n2094);
   U2566 : MUX2_X1 port map( A => REGISTERS_17_28_port, B => 
                           REGISTERS_18_28_port, S => n771, Z => n2095);
   U2567 : MUX2_X1 port map( A => REGISTERS_15_28_port, B => 
                           REGISTERS_16_28_port, S => n771, Z => n2096);
   U2568 : MUX2_X1 port map( A => n2096, B => n2095, S => n824, Z => n2097);
   U2569 : MUX2_X1 port map( A => n2097, B => n2094, S => n842, Z => n2098);
   U2570 : MUX2_X1 port map( A => n2098, B => n2091, S => n847, Z => n2099);
   U2571 : MUX2_X1 port map( A => REGISTERS_25_28_port, B => 
                           REGISTERS_26_28_port, S => n771, Z => n2100);
   U2572 : MUX2_X1 port map( A => REGISTERS_23_28_port, B => 
                           REGISTERS_24_28_port, S => n771, Z => n2101);
   U2573 : MUX2_X1 port map( A => n2101, B => n2100, S => n824, Z => n2102);
   U2574 : MUX2_X1 port map( A => REGISTERS_9_28_port, B => 
                           REGISTERS_10_28_port, S => n771, Z => n2103);
   U2575 : MUX2_X1 port map( A => REGISTERS_7_28_port, B => REGISTERS_8_28_port
                           , S => n771, Z => n2104);
   U2576 : MUX2_X1 port map( A => n2104, B => n2103, S => n825, Z => n2105);
   U2577 : MUX2_X1 port map( A => n2105, B => n2102, S => n842, Z => n2106);
   U2578 : MUX2_X1 port map( A => n2106, B => REGISTERS_39_28_port, S => n847, 
                           Z => n2107);
   U2579 : MUX2_X1 port map( A => n2107, B => n2099, S => n302, Z => n2108);
   U2580 : MUX2_X1 port map( A => n2108, B => n2089, S => n301, Z => N12233);
   U2581 : MUX2_X1 port map( A => REGISTERS_5_29_port, B => REGISTERS_6_29_port
                           , S => n771, Z => n2109);
   U2582 : MUX2_X1 port map( A => REGISTERS_3_29_port, B => REGISTERS_4_29_port
                           , S => n771, Z => n2110);
   U2583 : MUX2_X1 port map( A => n2110, B => n2109, S => n825, Z => n2111);
   U2584 : MUX2_X1 port map( A => REGISTERS_37_29_port, B => 
                           REGISTERS_38_29_port, S => n771, Z => n2112);
   U2585 : MUX2_X1 port map( A => REGISTERS_35_29_port, B => 
                           REGISTERS_36_29_port, S => n771, Z => n2113);
   U2586 : MUX2_X1 port map( A => n2113, B => n2112, S => n825, Z => n2114);
   U2587 : MUX2_X1 port map( A => REGISTERS_21_29_port, B => 
                           REGISTERS_22_29_port, S => n770, Z => n2115);
   U2588 : MUX2_X1 port map( A => REGISTERS_19_29_port, B => 
                           REGISTERS_20_29_port, S => n770, Z => n2116);
   U2589 : MUX2_X1 port map( A => n2116, B => n2115, S => n825, Z => n2117);
   U2590 : MUX2_X1 port map( A => n2117, B => n2114, S => n842, Z => n2118);
   U2591 : MUX2_X1 port map( A => n2118, B => n2111, S => n847, Z => n2119);
   U2592 : MUX2_X1 port map( A => REGISTERS_29_29_port, B => 
                           REGISTERS_30_29_port, S => n770, Z => n2120);
   U2593 : MUX2_X1 port map( A => REGISTERS_27_29_port, B => 
                           REGISTERS_28_29_port, S => n770, Z => n2121);
   U2594 : MUX2_X1 port map( A => n2121, B => n2120, S => n825, Z => n2122);
   U2595 : MUX2_X1 port map( A => REGISTERS_13_29_port, B => 
                           REGISTERS_14_29_port, S => n770, Z => n2123);
   U2596 : MUX2_X1 port map( A => REGISTERS_11_29_port, B => 
                           REGISTERS_12_29_port, S => n770, Z => n2124);
   U2597 : MUX2_X1 port map( A => n2124, B => n2123, S => n825, Z => n2125);
   U2598 : MUX2_X1 port map( A => n2125, B => n2122, S => n842, Z => n2126);
   U2599 : MUX2_X1 port map( A => n2126, B => n2119, S => n302, Z => n2127);
   U2600 : MUX2_X1 port map( A => REGISTERS_1_29_port, B => REGISTERS_2_29_port
                           , S => n770, Z => n2128);
   U2601 : MUX2_X1 port map( A => REGISTERS_0_29_port, B => n2128, S => n825, Z
                           => n2129);
   U2602 : MUX2_X1 port map( A => REGISTERS_33_29_port, B => 
                           REGISTERS_34_29_port, S => n770, Z => n2130);
   U2603 : MUX2_X1 port map( A => REGISTERS_31_29_port, B => 
                           REGISTERS_32_29_port, S => n770, Z => n2131);
   U2604 : MUX2_X1 port map( A => n2131, B => n2130, S => n825, Z => n2132);
   U2605 : MUX2_X1 port map( A => REGISTERS_17_29_port, B => 
                           REGISTERS_18_29_port, S => n770, Z => n2133);
   U2606 : MUX2_X1 port map( A => REGISTERS_15_29_port, B => 
                           REGISTERS_16_29_port, S => n770, Z => n2134);
   U2607 : MUX2_X1 port map( A => n2134, B => n2133, S => n825, Z => n2135);
   U2608 : MUX2_X1 port map( A => n2135, B => n2132, S => n842, Z => n2136);
   U2609 : MUX2_X1 port map( A => n2136, B => n2129, S => n847, Z => n2137);
   U2610 : MUX2_X1 port map( A => REGISTERS_25_29_port, B => 
                           REGISTERS_26_29_port, S => n770, Z => n2138);
   U2611 : MUX2_X1 port map( A => REGISTERS_23_29_port, B => 
                           REGISTERS_24_29_port, S => n769, Z => n2139);
   U2612 : MUX2_X1 port map( A => n2139, B => n2138, S => n825, Z => n2140);
   U2613 : MUX2_X1 port map( A => REGISTERS_9_29_port, B => 
                           REGISTERS_10_29_port, S => n769, Z => n2141);
   U2614 : MUX2_X1 port map( A => REGISTERS_7_29_port, B => REGISTERS_8_29_port
                           , S => n769, Z => n2142);
   U2615 : MUX2_X1 port map( A => n2142, B => n2141, S => n825, Z => n2143);
   U2616 : MUX2_X1 port map( A => n2143, B => n2140, S => n842, Z => n2144);
   U2617 : MUX2_X1 port map( A => n2144, B => REGISTERS_39_29_port, S => n847, 
                           Z => n2145);
   U2618 : MUX2_X1 port map( A => n2145, B => n2137, S => n302, Z => n2146);
   U2619 : MUX2_X1 port map( A => n2146, B => n2127, S => n301, Z => N12234);
   U2620 : MUX2_X1 port map( A => REGISTERS_5_30_port, B => REGISTERS_6_30_port
                           , S => n769, Z => n2147);
   U2621 : MUX2_X1 port map( A => REGISTERS_3_30_port, B => REGISTERS_4_30_port
                           , S => n769, Z => n2148);
   U2622 : MUX2_X1 port map( A => n2148, B => n2147, S => n825, Z => n2149);
   U2623 : MUX2_X1 port map( A => REGISTERS_37_30_port, B => 
                           REGISTERS_38_30_port, S => n769, Z => n2150);
   U2624 : MUX2_X1 port map( A => REGISTERS_35_30_port, B => 
                           REGISTERS_36_30_port, S => n769, Z => n2151);
   U2625 : MUX2_X1 port map( A => n2151, B => n2150, S => n826, Z => n2152);
   U2626 : MUX2_X1 port map( A => REGISTERS_21_30_port, B => 
                           REGISTERS_22_30_port, S => n769, Z => n2153);
   U2627 : MUX2_X1 port map( A => REGISTERS_19_30_port, B => 
                           REGISTERS_20_30_port, S => n769, Z => n2154);
   U2628 : MUX2_X1 port map( A => n2154, B => n2153, S => n826, Z => n2155);
   U2629 : MUX2_X1 port map( A => n2155, B => n2152, S => n842, Z => n2156);
   U2630 : MUX2_X1 port map( A => n2156, B => n2149, S => n847, Z => n2157);
   U2631 : MUX2_X1 port map( A => REGISTERS_29_30_port, B => 
                           REGISTERS_30_30_port, S => n769, Z => n2158);
   U2632 : MUX2_X1 port map( A => REGISTERS_27_30_port, B => 
                           REGISTERS_28_30_port, S => n769, Z => n2159);
   U2633 : MUX2_X1 port map( A => n2159, B => n2158, S => n826, Z => n2160);
   U2634 : MUX2_X1 port map( A => REGISTERS_13_30_port, B => 
                           REGISTERS_14_30_port, S => n769, Z => n2161);
   U2635 : MUX2_X1 port map( A => REGISTERS_11_30_port, B => 
                           REGISTERS_12_30_port, S => n768, Z => n2162);
   U2636 : MUX2_X1 port map( A => n2162, B => n2161, S => n826, Z => n2163);
   U2637 : MUX2_X1 port map( A => n2163, B => n2160, S => n842, Z => n2164);
   U2638 : MUX2_X1 port map( A => n2164, B => n2157, S => n302, Z => n2165);
   U2639 : MUX2_X1 port map( A => REGISTERS_1_30_port, B => REGISTERS_2_30_port
                           , S => n768, Z => n2166);
   U2640 : MUX2_X1 port map( A => REGISTERS_0_30_port, B => n2166, S => n826, Z
                           => n2167);
   U2641 : MUX2_X1 port map( A => REGISTERS_33_30_port, B => 
                           REGISTERS_34_30_port, S => n768, Z => n2168);
   U2642 : MUX2_X1 port map( A => REGISTERS_31_30_port, B => 
                           REGISTERS_32_30_port, S => n768, Z => n2169);
   U2643 : MUX2_X1 port map( A => n2169, B => n2168, S => n826, Z => n2170);
   U2644 : MUX2_X1 port map( A => REGISTERS_17_30_port, B => 
                           REGISTERS_18_30_port, S => n768, Z => n2171);
   U2645 : MUX2_X1 port map( A => REGISTERS_15_30_port, B => 
                           REGISTERS_16_30_port, S => n768, Z => n2172);
   U2646 : MUX2_X1 port map( A => n2172, B => n2171, S => n826, Z => n2173);
   U2647 : MUX2_X1 port map( A => n2173, B => n2170, S => n842, Z => n2174);
   U2648 : MUX2_X1 port map( A => n2174, B => n2167, S => n847, Z => n2175);
   U2649 : MUX2_X1 port map( A => REGISTERS_25_30_port, B => 
                           REGISTERS_26_30_port, S => n768, Z => n2176);
   U2650 : MUX2_X1 port map( A => REGISTERS_23_30_port, B => 
                           REGISTERS_24_30_port, S => n768, Z => n2177);
   U2651 : MUX2_X1 port map( A => n2177, B => n2176, S => n826, Z => n2178);
   U2652 : MUX2_X1 port map( A => REGISTERS_9_30_port, B => 
                           REGISTERS_10_30_port, S => n768, Z => n2179);
   U2653 : MUX2_X1 port map( A => REGISTERS_7_30_port, B => REGISTERS_8_30_port
                           , S => n768, Z => n2180);
   U2654 : MUX2_X1 port map( A => n2180, B => n2179, S => n826, Z => n2181);
   U2655 : MUX2_X1 port map( A => n2181, B => n2178, S => n842, Z => n2182);
   U2656 : MUX2_X1 port map( A => n2182, B => REGISTERS_39_30_port, S => n847, 
                           Z => n2183);
   U2657 : MUX2_X1 port map( A => n2183, B => n2175, S => n302, Z => n2184);
   U2658 : MUX2_X1 port map( A => n2184, B => n2165, S => n301, Z => N12235);
   U2659 : MUX2_X1 port map( A => REGISTERS_5_31_port, B => REGISTERS_6_31_port
                           , S => n768, Z => n2185);
   U2660 : MUX2_X1 port map( A => REGISTERS_3_31_port, B => REGISTERS_4_31_port
                           , S => n768, Z => n2186);
   U2661 : MUX2_X1 port map( A => n2186, B => n2185, S => n826, Z => n2187);
   U2662 : MUX2_X1 port map( A => REGISTERS_37_31_port, B => 
                           REGISTERS_38_31_port, S => n767, Z => n2188);
   U2663 : MUX2_X1 port map( A => REGISTERS_35_31_port, B => 
                           REGISTERS_36_31_port, S => n767, Z => n2189);
   U2664 : MUX2_X1 port map( A => n2189, B => n2188, S => n826, Z => n2190);
   U2665 : MUX2_X1 port map( A => REGISTERS_21_31_port, B => 
                           REGISTERS_22_31_port, S => n767, Z => n2191);
   U2666 : MUX2_X1 port map( A => REGISTERS_19_31_port, B => 
                           REGISTERS_20_31_port, S => n767, Z => n2192);
   U2667 : MUX2_X1 port map( A => n2192, B => n2191, S => n826, Z => n2193);
   U2668 : MUX2_X1 port map( A => n2193, B => n2190, S => n842, Z => n2194);
   U2669 : MUX2_X1 port map( A => n2194, B => n2187, S => n847, Z => n2195);
   U2670 : MUX2_X1 port map( A => REGISTERS_29_31_port, B => 
                           REGISTERS_30_31_port, S => n767, Z => n2196);
   U2671 : MUX2_X1 port map( A => REGISTERS_27_31_port, B => 
                           REGISTERS_28_31_port, S => n767, Z => n2197);
   U2672 : MUX2_X1 port map( A => n2197, B => n2196, S => n827, Z => n2198);
   U2673 : MUX2_X1 port map( A => REGISTERS_13_31_port, B => 
                           REGISTERS_14_31_port, S => n767, Z => n2199);
   U2674 : MUX2_X1 port map( A => REGISTERS_11_31_port, B => 
                           REGISTERS_12_31_port, S => n767, Z => n2200);
   U2675 : MUX2_X1 port map( A => n2200, B => n2199, S => n827, Z => n2201);
   U2676 : MUX2_X1 port map( A => n2201, B => n2198, S => n842, Z => n2202);
   U2677 : MUX2_X1 port map( A => n2202, B => n2195, S => n302, Z => n2203);
   U2678 : MUX2_X1 port map( A => REGISTERS_1_31_port, B => REGISTERS_2_31_port
                           , S => n767, Z => n2204);
   U2679 : MUX2_X1 port map( A => REGISTERS_0_31_port, B => n2204, S => n827, Z
                           => n2205);
   U2680 : MUX2_X1 port map( A => REGISTERS_33_31_port, B => 
                           REGISTERS_34_31_port, S => n767, Z => n2206);
   U2681 : MUX2_X1 port map( A => REGISTERS_31_31_port, B => 
                           REGISTERS_32_31_port, S => n767, Z => n2207);
   U2682 : MUX2_X1 port map( A => n2207, B => n2206, S => n827, Z => n2208);
   U2683 : MUX2_X1 port map( A => REGISTERS_17_31_port, B => 
                           REGISTERS_18_31_port, S => n767, Z => n2209);
   U2684 : MUX2_X1 port map( A => REGISTERS_15_31_port, B => 
                           REGISTERS_16_31_port, S => n766, Z => n2210);
   U2685 : MUX2_X1 port map( A => n2210, B => n2209, S => n827, Z => n2211);
   U2686 : MUX2_X1 port map( A => n2211, B => n2208, S => n842, Z => n2212);
   U2687 : MUX2_X1 port map( A => n2212, B => n2205, S => n847, Z => n2213);
   U2688 : MUX2_X1 port map( A => REGISTERS_25_31_port, B => 
                           REGISTERS_26_31_port, S => n766, Z => n2214);
   U2689 : MUX2_X1 port map( A => REGISTERS_23_31_port, B => 
                           REGISTERS_24_31_port, S => n773, Z => n2215);
   U2690 : MUX2_X1 port map( A => n2215, B => n2214, S => n814, Z => n2216);
   U2691 : MUX2_X1 port map( A => REGISTERS_9_31_port, B => 
                           REGISTERS_10_31_port, S => n754, Z => n2217);
   U2692 : MUX2_X1 port map( A => REGISTERS_7_31_port, B => REGISTERS_8_31_port
                           , S => n779, Z => n2218);
   U2693 : MUX2_X1 port map( A => n2218, B => n2217, S => n827, Z => n2219);
   U2694 : MUX2_X1 port map( A => n2219, B => n2216, S => n841, Z => n2220);
   U2695 : MUX2_X1 port map( A => n2220, B => REGISTERS_39_31_port, S => n846, 
                           Z => n2221);
   U2696 : MUX2_X1 port map( A => n2221, B => n2213, S => n302, Z => n2222);
   U2697 : MUX2_X1 port map( A => n2222, B => n2203, S => n301, Z => N12236);
   U2698 : MUX2_X1 port map( A => n1038, B => REGISTERS_39_0_port, S => n841, Z
                           => n2223);
   U2699 : MUX2_X1 port map( A => n2223, B => n1041, S => n846, Z => n2224);
   U2700 : MUX2_X1 port map( A => n1035, B => n2224, S => n302, Z => n2225);
   U2701 : MUX2_X1 port map( A => n1025, B => n2225, S => n301, Z => N5250);
   U2702 : MUX2_X1 port map( A => n1076, B => REGISTERS_39_1_port, S => n841, Z
                           => n2226);
   U2703 : MUX2_X1 port map( A => n2226, B => n1079, S => n846, Z => n2227);
   U2704 : MUX2_X1 port map( A => n1073, B => n2227, S => n302, Z => n2228);
   U2705 : MUX2_X1 port map( A => n1063, B => n2228, S => n301, Z => N5251);
   U2706 : MUX2_X1 port map( A => n1114, B => REGISTERS_39_2_port, S => n841, Z
                           => n2229);
   U2707 : MUX2_X1 port map( A => n2229, B => n1117, S => n846, Z => n2230);
   U2708 : MUX2_X1 port map( A => n1111, B => n2230, S => n302, Z => n2231);
   U2709 : MUX2_X1 port map( A => n1101, B => n2231, S => n301, Z => N5252);
   U2710 : MUX2_X1 port map( A => n1152, B => REGISTERS_39_3_port, S => n841, Z
                           => n2232);
   U2711 : MUX2_X1 port map( A => n2232, B => n1155, S => n846, Z => n2233);
   U2712 : MUX2_X1 port map( A => n1149, B => n2233, S => n302, Z => n2234);
   U2713 : MUX2_X1 port map( A => n1139, B => n2234, S => n301, Z => N5253);
   U2714 : MUX2_X1 port map( A => n1190, B => REGISTERS_39_4_port, S => n841, Z
                           => n2235);
   U2715 : MUX2_X1 port map( A => n2235, B => n1193, S => n846, Z => n2236);
   U2716 : MUX2_X1 port map( A => n1187, B => n2236, S => n302, Z => n2237);
   U2717 : MUX2_X1 port map( A => n1177, B => n2237, S => n301, Z => N5254);
   U2718 : MUX2_X1 port map( A => n1228, B => REGISTERS_39_5_port, S => n841, Z
                           => n2238);
   U2719 : MUX2_X1 port map( A => n2238, B => n1231, S => n846, Z => n2239);
   U2720 : MUX2_X1 port map( A => n1225, B => n2239, S => n302, Z => n2240);
   U2721 : MUX2_X1 port map( A => n1215, B => n2240, S => n301, Z => N5255);
   U2722 : MUX2_X1 port map( A => n1266, B => REGISTERS_39_6_port, S => n841, Z
                           => n2241);
   U2723 : MUX2_X1 port map( A => n2241, B => n1269, S => n846, Z => n2242);
   U2724 : MUX2_X1 port map( A => n1263, B => n2242, S => n302, Z => n2243);
   U2725 : MUX2_X1 port map( A => n1253, B => n2243, S => n301, Z => N5256);
   U2726 : MUX2_X1 port map( A => n1304, B => REGISTERS_39_7_port, S => n841, Z
                           => n2244);
   U2727 : MUX2_X1 port map( A => n2244, B => n1307, S => n846, Z => n2245);
   U2728 : MUX2_X1 port map( A => n1301, B => n2245, S => n302, Z => n2246);
   U2729 : MUX2_X1 port map( A => n1291, B => n2246, S => n301, Z => N5257);
   U2730 : MUX2_X1 port map( A => n1342, B => REGISTERS_39_8_port, S => n841, Z
                           => n2247);
   U2731 : MUX2_X1 port map( A => n2247, B => n1345, S => n846, Z => n2248);
   U2732 : MUX2_X1 port map( A => n1339, B => n2248, S => n302, Z => n2249);
   U2733 : MUX2_X1 port map( A => n1329, B => n2249, S => n301, Z => N5258);
   U2734 : MUX2_X1 port map( A => n1380, B => REGISTERS_39_9_port, S => n841, Z
                           => n2250);
   U2735 : MUX2_X1 port map( A => n2250, B => n1383, S => n846, Z => n2251);
   U2736 : MUX2_X1 port map( A => n1377, B => n2251, S => n302, Z => n2252);
   U2737 : MUX2_X1 port map( A => n1367, B => n2252, S => n301, Z => N5259);
   U2738 : MUX2_X1 port map( A => n1418, B => REGISTERS_39_10_port, S => n841, 
                           Z => n2253);
   U2739 : MUX2_X1 port map( A => n2253, B => n1421, S => n846, Z => n2254);
   U2740 : MUX2_X1 port map( A => n1415, B => n2254, S => n302, Z => n2255);
   U2741 : MUX2_X1 port map( A => n1405, B => n2255, S => n301, Z => N5260);
   U2742 : MUX2_X1 port map( A => n1456, B => REGISTERS_39_11_port, S => n841, 
                           Z => n2256);
   U2743 : MUX2_X1 port map( A => n2256, B => n1459, S => n846, Z => n2257);
   U2744 : MUX2_X1 port map( A => n1453, B => n2257, S => n302, Z => n2258);
   U2745 : MUX2_X1 port map( A => n1443, B => n2258, S => n301, Z => N5261);
   U2746 : MUX2_X1 port map( A => n1494, B => REGISTERS_39_12_port, S => n841, 
                           Z => n2259);
   U2747 : MUX2_X1 port map( A => n2259, B => n1497, S => n846, Z => n2260);
   U2748 : MUX2_X1 port map( A => n1491, B => n2260, S => n302, Z => n2261);
   U2749 : MUX2_X1 port map( A => n1481, B => n2261, S => n301, Z => N5262);
   U2750 : MUX2_X1 port map( A => n1532, B => REGISTERS_39_13_port, S => n841, 
                           Z => n2262);
   U2751 : MUX2_X1 port map( A => n2262, B => n1535, S => n846, Z => n2263);
   U2752 : MUX2_X1 port map( A => n1529, B => n2263, S => n302, Z => n2264);
   U2753 : MUX2_X1 port map( A => n1519, B => n2264, S => n301, Z => N5263);
   U2754 : MUX2_X1 port map( A => n1570, B => REGISTERS_39_14_port, S => n841, 
                           Z => n2265);
   U2755 : MUX2_X1 port map( A => n2265, B => n1573, S => n846, Z => n2266);
   U2756 : MUX2_X1 port map( A => n1567, B => n2266, S => n302, Z => n2267);
   U2757 : MUX2_X1 port map( A => n1557, B => n2267, S => n301, Z => N5264);
   U2758 : MUX2_X1 port map( A => n1608, B => REGISTERS_39_15_port, S => n841, 
                           Z => n2268);
   U2759 : MUX2_X1 port map( A => n2268, B => n1611, S => n846, Z => n2269);
   U2760 : MUX2_X1 port map( A => n1605, B => n2269, S => n302, Z => n2270);
   U2761 : MUX2_X1 port map( A => n1595, B => n2270, S => n301, Z => N5265);
   U2762 : MUX2_X1 port map( A => n1646, B => REGISTERS_39_16_port, S => n841, 
                           Z => n2271);
   U2763 : MUX2_X1 port map( A => n2271, B => n1649, S => n846, Z => n2272);
   U2764 : MUX2_X1 port map( A => n1643, B => n2272, S => n302, Z => n2273);
   U2765 : MUX2_X1 port map( A => n1633, B => n2273, S => n301, Z => N5266);
   U2766 : MUX2_X1 port map( A => n1684, B => REGISTERS_39_17_port, S => n841, 
                           Z => n2274);
   U2767 : MUX2_X1 port map( A => n2274, B => n1687, S => n846, Z => n2275);
   U2768 : MUX2_X1 port map( A => n1681, B => n2275, S => n302, Z => n2276);
   U2769 : MUX2_X1 port map( A => n1671, B => n2276, S => n301, Z => N5267);
   U2770 : MUX2_X1 port map( A => n1722, B => REGISTERS_39_18_port, S => n841, 
                           Z => n2277);
   U2771 : MUX2_X1 port map( A => n2277, B => n1725, S => n846, Z => n2278);
   U2772 : MUX2_X1 port map( A => n1719, B => n2278, S => n302, Z => n2279);
   U2773 : MUX2_X1 port map( A => n1709, B => n2279, S => n301, Z => N5268);
   U2774 : MUX2_X1 port map( A => n1760, B => REGISTERS_39_19_port, S => n841, 
                           Z => n2280);
   U2775 : MUX2_X1 port map( A => n2280, B => n1763, S => n846, Z => n2281);
   U2776 : MUX2_X1 port map( A => n1757, B => n2281, S => n302, Z => n2282);
   U2777 : MUX2_X1 port map( A => n1747, B => n2282, S => n301, Z => N5269);
   U2778 : MUX2_X1 port map( A => n1798, B => REGISTERS_39_20_port, S => n841, 
                           Z => n2283);
   U2779 : MUX2_X1 port map( A => n2283, B => n1801, S => n846, Z => n2284);
   U2780 : MUX2_X1 port map( A => n1795, B => n2284, S => n302, Z => n2285);
   U2781 : MUX2_X1 port map( A => n1785, B => n2285, S => n301, Z => N5270);
   U2782 : MUX2_X1 port map( A => n1836, B => REGISTERS_39_21_port, S => n841, 
                           Z => n2286);
   U2783 : MUX2_X1 port map( A => n2286, B => n1839, S => n846, Z => n2287);
   U2784 : MUX2_X1 port map( A => n1833, B => n2287, S => n302, Z => n2288);
   U2785 : MUX2_X1 port map( A => n1823, B => n2288, S => n301, Z => N5271);
   U2786 : MUX2_X1 port map( A => n1874, B => REGISTERS_39_22_port, S => n841, 
                           Z => n2289);
   U2787 : MUX2_X1 port map( A => n2289, B => n1877, S => n846, Z => n2290);
   U2788 : MUX2_X1 port map( A => n1871, B => n2290, S => n302, Z => n2291);
   U2789 : MUX2_X1 port map( A => n1861, B => n2291, S => n301, Z => N5272);
   U2790 : MUX2_X1 port map( A => n1912, B => REGISTERS_39_23_port, S => n841, 
                           Z => n2292);
   U2791 : MUX2_X1 port map( A => n2292, B => n1915, S => n846, Z => n2293);
   U2792 : MUX2_X1 port map( A => n1909, B => n2293, S => n302, Z => n2294);
   U2793 : MUX2_X1 port map( A => n1899, B => n2294, S => n301, Z => N5273);
   U2794 : MUX2_X1 port map( A => n1950, B => REGISTERS_39_24_port, S => n841, 
                           Z => n2295);
   U2795 : MUX2_X1 port map( A => n2295, B => n1953, S => n846, Z => n2296);
   U2796 : MUX2_X1 port map( A => n1947, B => n2296, S => n302, Z => n2297);
   U2797 : MUX2_X1 port map( A => n1937, B => n2297, S => n301, Z => N5274);
   U2798 : MUX2_X1 port map( A => n1988, B => REGISTERS_39_25_port, S => n841, 
                           Z => n2298);
   U2799 : MUX2_X1 port map( A => n2298, B => n1991, S => n846, Z => n2299);
   U2800 : MUX2_X1 port map( A => n1985, B => n2299, S => n302, Z => n2300);
   U2801 : MUX2_X1 port map( A => n1975, B => n2300, S => n301, Z => N5275);
   U2802 : MUX2_X1 port map( A => n2026, B => REGISTERS_39_26_port, S => n841, 
                           Z => n2301);
   U2803 : MUX2_X1 port map( A => n2301, B => n2029, S => n846, Z => n2302);
   U2804 : MUX2_X1 port map( A => n2023, B => n2302, S => n302, Z => n2303);
   U2805 : MUX2_X1 port map( A => n2013, B => n2303, S => n301, Z => N5276);
   U2806 : MUX2_X1 port map( A => n2064, B => REGISTERS_39_27_port, S => n841, 
                           Z => n2304);
   U2807 : MUX2_X1 port map( A => n2304, B => n2067, S => n846, Z => n2305);
   U2808 : MUX2_X1 port map( A => n2061, B => n2305, S => n302, Z => n2306);
   U2809 : MUX2_X1 port map( A => n2051, B => n2306, S => n301, Z => N5277);
   U2810 : MUX2_X1 port map( A => n2102, B => REGISTERS_39_28_port, S => n841, 
                           Z => n2307);
   U2811 : MUX2_X1 port map( A => n2307, B => n2105, S => n846, Z => n2308);
   U2812 : MUX2_X1 port map( A => n2099, B => n2308, S => n302, Z => n2309);
   U2813 : MUX2_X1 port map( A => n2089, B => n2309, S => n301, Z => N5278);
   U2814 : MUX2_X1 port map( A => n2140, B => REGISTERS_39_29_port, S => n841, 
                           Z => n2310);
   U2815 : MUX2_X1 port map( A => n2310, B => n2143, S => n846, Z => n2311);
   U2816 : MUX2_X1 port map( A => n2137, B => n2311, S => n302, Z => n2312);
   U2817 : MUX2_X1 port map( A => n2127, B => n2312, S => n301, Z => N5279);
   U2818 : MUX2_X1 port map( A => n2178, B => REGISTERS_39_30_port, S => n841, 
                           Z => n2313);
   U2819 : MUX2_X1 port map( A => n2313, B => n2181, S => n846, Z => n2314);
   U2820 : MUX2_X1 port map( A => n2175, B => n2314, S => n302, Z => n2315);
   U2821 : MUX2_X1 port map( A => n2165, B => n2315, S => n301, Z => N5280);
   U2822 : MUX2_X1 port map( A => n2216, B => REGISTERS_39_31_port, S => n843, 
                           Z => n2316);
   U2823 : MUX2_X1 port map( A => n2316, B => n2219, S => n847, Z => n2317);
   U2824 : MUX2_X1 port map( A => n2213, B => n2317, S => n302, Z => n2318);
   U2825 : MUX2_X1 port map( A => n2203, B => n2318, S => n301, Z => N5281);
   U2826 : MUX2_X1 port map( A => REGISTERS_37_0_port, B => REGISTERS_39_0_port
                           , S => n636, Z => n2319);
   U2827 : MUX2_X1 port map( A => REGISTERS_36_0_port, B => REGISTERS_38_0_port
                           , S => n636, Z => n2320);
   U2828 : MUX2_X1 port map( A => n2320, B => n2319, S => n667, Z => n2321);
   U2829 : MUX2_X1 port map( A => REGISTERS_33_0_port, B => REGISTERS_35_0_port
                           , S => n636, Z => n2322);
   U2830 : MUX2_X1 port map( A => REGISTERS_32_0_port, B => REGISTERS_34_0_port
                           , S => n636, Z => n2323);
   U2831 : MUX2_X1 port map( A => n2323, B => n2322, S => n667, Z => n2324);
   U2832 : MUX2_X1 port map( A => n2324, B => n2321, S => n593, Z => n2325);
   U2833 : MUX2_X1 port map( A => REGISTERS_29_0_port, B => REGISTERS_31_0_port
                           , S => n636, Z => n2326);
   U2834 : MUX2_X1 port map( A => REGISTERS_28_0_port, B => REGISTERS_30_0_port
                           , S => n636, Z => n2327);
   U2835 : MUX2_X1 port map( A => n2327, B => n2326, S => n667, Z => n2328);
   U2836 : MUX2_X1 port map( A => REGISTERS_25_0_port, B => REGISTERS_27_0_port
                           , S => n636, Z => n2329);
   U2837 : MUX2_X1 port map( A => REGISTERS_24_0_port, B => REGISTERS_26_0_port
                           , S => n636, Z => n2330);
   U2838 : MUX2_X1 port map( A => n2330, B => n2329, S => n667, Z => n2331);
   U2839 : MUX2_X1 port map( A => n2331, B => n2328, S => n593, Z => n2332);
   U2840 : MUX2_X1 port map( A => REGISTERS_21_0_port, B => REGISTERS_23_0_port
                           , S => n636, Z => n2333);
   U2841 : MUX2_X1 port map( A => REGISTERS_20_0_port, B => REGISTERS_22_0_port
                           , S => n636, Z => n2334);
   U2842 : MUX2_X1 port map( A => n2334, B => n2333, S => n667, Z => n2335);
   U2843 : MUX2_X1 port map( A => REGISTERS_17_0_port, B => REGISTERS_19_0_port
                           , S => n636, Z => n2336);
   U2844 : MUX2_X1 port map( A => REGISTERS_16_0_port, B => REGISTERS_18_0_port
                           , S => n636, Z => n2337);
   U2845 : MUX2_X1 port map( A => n2337, B => n2336, S => n667, Z => n2338);
   U2846 : MUX2_X1 port map( A => n2338, B => n2335, S => n593, Z => n2339);
   U2847 : MUX2_X1 port map( A => n2339, B => n2332, S => r3013_A_3_port, Z => 
                           n2340);
   U2848 : MUX2_X1 port map( A => REGISTERS_13_0_port, B => REGISTERS_15_0_port
                           , S => n635, Z => n2341);
   U2849 : MUX2_X1 port map( A => REGISTERS_12_0_port, B => REGISTERS_14_0_port
                           , S => n635, Z => n2342);
   U2850 : MUX2_X1 port map( A => n2342, B => n2341, S => n667, Z => n2343);
   U2851 : MUX2_X1 port map( A => REGISTERS_9_0_port, B => REGISTERS_11_0_port,
                           S => n635, Z => n2344);
   U2852 : MUX2_X1 port map( A => REGISTERS_8_0_port, B => REGISTERS_10_0_port,
                           S => n635, Z => n2345);
   U2853 : MUX2_X1 port map( A => n2345, B => n2344, S => n666, Z => n2346);
   U2854 : MUX2_X1 port map( A => n2346, B => n2343, S => n593, Z => n2347);
   U2855 : MUX2_X1 port map( A => REGISTERS_5_0_port, B => REGISTERS_7_0_port, 
                           S => n635, Z => n2348);
   U2856 : MUX2_X1 port map( A => REGISTERS_4_0_port, B => REGISTERS_6_0_port, 
                           S => n635, Z => n2349);
   U2857 : MUX2_X1 port map( A => n2349, B => n2348, S => n666, Z => n2350);
   U2858 : MUX2_X1 port map( A => REGISTERS_1_0_port, B => REGISTERS_3_0_port, 
                           S => n635, Z => n2351);
   U2859 : MUX2_X1 port map( A => REGISTERS_0_0_port, B => REGISTERS_2_0_port, 
                           S => n635, Z => n2352);
   U2860 : MUX2_X1 port map( A => n2352, B => n2351, S => n666, Z => n2353);
   U2861 : MUX2_X1 port map( A => n2353, B => n2350, S => n593, Z => n2354);
   U2862 : MUX2_X1 port map( A => n2354, B => n2347, S => r3013_A_3_port, Z => 
                           n2355);
   U2863 : MUX2_X1 port map( A => n2355, B => n2340, S => r3013_A_4_port, Z => 
                           n2356);
   U2864 : MUX2_X1 port map( A => n2356, B => n2325, S => ADD_RD2_5_port, Z => 
                           N4526);
   U2865 : MUX2_X1 port map( A => REGISTERS_37_1_port, B => REGISTERS_39_1_port
                           , S => n635, Z => n2357);
   U2866 : MUX2_X1 port map( A => REGISTERS_36_1_port, B => REGISTERS_38_1_port
                           , S => n635, Z => n2358);
   U2867 : MUX2_X1 port map( A => n2358, B => n2357, S => n666, Z => n2359);
   U2868 : MUX2_X1 port map( A => REGISTERS_33_1_port, B => REGISTERS_35_1_port
                           , S => n635, Z => n2360);
   U2869 : MUX2_X1 port map( A => REGISTERS_32_1_port, B => REGISTERS_34_1_port
                           , S => n635, Z => n2361);
   U2870 : MUX2_X1 port map( A => n2361, B => n2360, S => n666, Z => n2362);
   U2871 : MUX2_X1 port map( A => n2362, B => n2359, S => n592, Z => n2363);
   U2872 : MUX2_X1 port map( A => REGISTERS_29_1_port, B => REGISTERS_31_1_port
                           , S => n635, Z => n2364);
   U2873 : MUX2_X1 port map( A => REGISTERS_28_1_port, B => REGISTERS_30_1_port
                           , S => n635, Z => n2365);
   U2874 : MUX2_X1 port map( A => n2365, B => n2364, S => n666, Z => n2366);
   U2875 : MUX2_X1 port map( A => REGISTERS_25_1_port, B => REGISTERS_27_1_port
                           , S => n635, Z => n2367);
   U2876 : MUX2_X1 port map( A => REGISTERS_24_1_port, B => REGISTERS_26_1_port
                           , S => n634, Z => n2368);
   U2877 : MUX2_X1 port map( A => n2368, B => n2367, S => n666, Z => n2369);
   U2878 : MUX2_X1 port map( A => n2369, B => n2366, S => n592, Z => n2370);
   U2879 : MUX2_X1 port map( A => REGISTERS_21_1_port, B => REGISTERS_23_1_port
                           , S => n634, Z => n2371);
   U2880 : MUX2_X1 port map( A => REGISTERS_20_1_port, B => REGISTERS_22_1_port
                           , S => n634, Z => n2372);
   U2881 : MUX2_X1 port map( A => n2372, B => n2371, S => n666, Z => n2373);
   U2882 : MUX2_X1 port map( A => REGISTERS_17_1_port, B => REGISTERS_19_1_port
                           , S => n634, Z => n2374);
   U2883 : MUX2_X1 port map( A => REGISTERS_16_1_port, B => REGISTERS_18_1_port
                           , S => n634, Z => n2375);
   U2884 : MUX2_X1 port map( A => n2375, B => n2374, S => n666, Z => n2376);
   U2885 : MUX2_X1 port map( A => n2376, B => n2373, S => n592, Z => n2377);
   U2886 : MUX2_X1 port map( A => n2377, B => n2370, S => r3013_A_3_port, Z => 
                           n2378);
   U2887 : MUX2_X1 port map( A => REGISTERS_13_1_port, B => REGISTERS_15_1_port
                           , S => n634, Z => n2379);
   U2888 : MUX2_X1 port map( A => REGISTERS_12_1_port, B => REGISTERS_14_1_port
                           , S => n634, Z => n2380);
   U2889 : MUX2_X1 port map( A => n2380, B => n2379, S => n666, Z => n2381);
   U2890 : MUX2_X1 port map( A => REGISTERS_9_1_port, B => REGISTERS_11_1_port,
                           S => n634, Z => n2382);
   U2891 : MUX2_X1 port map( A => REGISTERS_8_1_port, B => REGISTERS_10_1_port,
                           S => n634, Z => n2383);
   U2892 : MUX2_X1 port map( A => n2383, B => n2382, S => n666, Z => n2384);
   U2893 : MUX2_X1 port map( A => n2384, B => n2381, S => n592, Z => n2385);
   U2894 : MUX2_X1 port map( A => REGISTERS_5_1_port, B => REGISTERS_7_1_port, 
                           S => n634, Z => n2386);
   U2895 : MUX2_X1 port map( A => REGISTERS_4_1_port, B => REGISTERS_6_1_port, 
                           S => n634, Z => n2387);
   U2896 : MUX2_X1 port map( A => n2387, B => n2386, S => n666, Z => n2388);
   U2897 : MUX2_X1 port map( A => REGISTERS_1_1_port, B => REGISTERS_3_1_port, 
                           S => n634, Z => n2389);
   U2898 : MUX2_X1 port map( A => REGISTERS_0_1_port, B => REGISTERS_2_1_port, 
                           S => n634, Z => n2390);
   U2899 : MUX2_X1 port map( A => n2390, B => n2389, S => n666, Z => n2391);
   U2900 : MUX2_X1 port map( A => n2391, B => n2388, S => n592, Z => n2392);
   U2901 : MUX2_X1 port map( A => n2392, B => n2385, S => r3013_A_3_port, Z => 
                           n2393);
   U2902 : MUX2_X1 port map( A => n2393, B => n2378, S => r3013_A_4_port, Z => 
                           n2394);
   U2903 : MUX2_X1 port map( A => n2394, B => n2363, S => ADD_RD2_5_port, Z => 
                           N4525);
   U2904 : MUX2_X1 port map( A => REGISTERS_37_2_port, B => REGISTERS_39_2_port
                           , S => n634, Z => n2395);
   U2905 : MUX2_X1 port map( A => REGISTERS_36_2_port, B => REGISTERS_38_2_port
                           , S => n634, Z => n2396);
   U2906 : MUX2_X1 port map( A => n2396, B => n2395, S => n666, Z => n2397);
   U2907 : MUX2_X1 port map( A => REGISTERS_33_2_port, B => REGISTERS_35_2_port
                           , S => n633, Z => n2398);
   U2908 : MUX2_X1 port map( A => REGISTERS_32_2_port, B => REGISTERS_34_2_port
                           , S => n633, Z => n2399);
   U2909 : MUX2_X1 port map( A => n2399, B => n2398, S => n666, Z => n2400);
   U2910 : MUX2_X1 port map( A => n2400, B => n2397, S => n592, Z => n2401);
   U2911 : MUX2_X1 port map( A => REGISTERS_29_2_port, B => REGISTERS_31_2_port
                           , S => n633, Z => n2402);
   U2912 : MUX2_X1 port map( A => REGISTERS_28_2_port, B => REGISTERS_30_2_port
                           , S => n633, Z => n2403);
   U2913 : MUX2_X1 port map( A => n2403, B => n2402, S => n665, Z => n2404);
   U2914 : MUX2_X1 port map( A => REGISTERS_25_2_port, B => REGISTERS_27_2_port
                           , S => n633, Z => n2405);
   U2915 : MUX2_X1 port map( A => REGISTERS_24_2_port, B => REGISTERS_26_2_port
                           , S => n633, Z => n2406);
   U2916 : MUX2_X1 port map( A => n2406, B => n2405, S => n665, Z => n2407);
   U2917 : MUX2_X1 port map( A => n2407, B => n2404, S => n592, Z => n2408);
   U2918 : MUX2_X1 port map( A => REGISTERS_21_2_port, B => REGISTERS_23_2_port
                           , S => n633, Z => n2409);
   U2919 : MUX2_X1 port map( A => REGISTERS_20_2_port, B => REGISTERS_22_2_port
                           , S => n633, Z => n2410);
   U2920 : MUX2_X1 port map( A => n2410, B => n2409, S => n665, Z => n2411);
   U2921 : MUX2_X1 port map( A => REGISTERS_17_2_port, B => REGISTERS_19_2_port
                           , S => n633, Z => n2412);
   U2922 : MUX2_X1 port map( A => REGISTERS_16_2_port, B => REGISTERS_18_2_port
                           , S => n633, Z => n2413);
   U2923 : MUX2_X1 port map( A => n2413, B => n2412, S => n665, Z => n2414);
   U2924 : MUX2_X1 port map( A => n2414, B => n2411, S => n592, Z => n2415);
   U2925 : MUX2_X1 port map( A => n2415, B => n2408, S => r3013_A_3_port, Z => 
                           n2416);
   U2926 : MUX2_X1 port map( A => REGISTERS_13_2_port, B => REGISTERS_15_2_port
                           , S => n633, Z => n2417);
   U2927 : MUX2_X1 port map( A => REGISTERS_12_2_port, B => REGISTERS_14_2_port
                           , S => n633, Z => n2418);
   U2928 : MUX2_X1 port map( A => n2418, B => n2417, S => n665, Z => n2419);
   U2929 : MUX2_X1 port map( A => REGISTERS_9_2_port, B => REGISTERS_11_2_port,
                           S => n633, Z => n2420);
   U2930 : MUX2_X1 port map( A => REGISTERS_8_2_port, B => REGISTERS_10_2_port,
                           S => n633, Z => n2421);
   U2931 : MUX2_X1 port map( A => n2421, B => n2420, S => n665, Z => n2422);
   U2932 : MUX2_X1 port map( A => n2422, B => n2419, S => n592, Z => n2423);
   U2933 : MUX2_X1 port map( A => REGISTERS_5_2_port, B => REGISTERS_7_2_port, 
                           S => n633, Z => n2424);
   U2934 : MUX2_X1 port map( A => REGISTERS_4_2_port, B => REGISTERS_6_2_port, 
                           S => n632, Z => n2425);
   U2935 : MUX2_X1 port map( A => n2425, B => n2424, S => n665, Z => n2426);
   U2936 : MUX2_X1 port map( A => REGISTERS_1_2_port, B => REGISTERS_3_2_port, 
                           S => n632, Z => n2427);
   U2937 : MUX2_X1 port map( A => REGISTERS_0_2_port, B => REGISTERS_2_2_port, 
                           S => n632, Z => n2428);
   U2938 : MUX2_X1 port map( A => n2428, B => n2427, S => n665, Z => n2429);
   U2939 : MUX2_X1 port map( A => n2429, B => n2426, S => n592, Z => n2430);
   U2940 : MUX2_X1 port map( A => n2430, B => n2423, S => r3013_A_3_port, Z => 
                           n2431);
   U2941 : MUX2_X1 port map( A => n2431, B => n2416, S => r3013_A_4_port, Z => 
                           n2432);
   U2942 : MUX2_X1 port map( A => n2432, B => n2401, S => ADD_RD2_5_port, Z => 
                           N4524);
   U2943 : MUX2_X1 port map( A => REGISTERS_37_3_port, B => REGISTERS_39_3_port
                           , S => n632, Z => n2433);
   U2944 : MUX2_X1 port map( A => REGISTERS_36_3_port, B => REGISTERS_38_3_port
                           , S => n632, Z => n2434);
   U2945 : MUX2_X1 port map( A => n2434, B => n2433, S => n665, Z => n2435);
   U2946 : MUX2_X1 port map( A => REGISTERS_33_3_port, B => REGISTERS_35_3_port
                           , S => n632, Z => n2436);
   U2947 : MUX2_X1 port map( A => REGISTERS_32_3_port, B => REGISTERS_34_3_port
                           , S => n632, Z => n2437);
   U2948 : MUX2_X1 port map( A => n2437, B => n2436, S => n665, Z => n2438);
   U2949 : MUX2_X1 port map( A => n2438, B => n2435, S => n592, Z => n2439);
   U2950 : MUX2_X1 port map( A => REGISTERS_29_3_port, B => REGISTERS_31_3_port
                           , S => n632, Z => n2440);
   U2951 : MUX2_X1 port map( A => REGISTERS_28_3_port, B => REGISTERS_30_3_port
                           , S => n632, Z => n2441);
   U2952 : MUX2_X1 port map( A => n2441, B => n2440, S => n665, Z => n2442);
   U2953 : MUX2_X1 port map( A => REGISTERS_25_3_port, B => REGISTERS_27_3_port
                           , S => n632, Z => n2443);
   U2954 : MUX2_X1 port map( A => REGISTERS_24_3_port, B => REGISTERS_26_3_port
                           , S => n632, Z => n2444);
   U2955 : MUX2_X1 port map( A => n2444, B => n2443, S => n665, Z => n2445);
   U2956 : MUX2_X1 port map( A => n2445, B => n2442, S => n592, Z => n2446);
   U2957 : MUX2_X1 port map( A => REGISTERS_21_3_port, B => REGISTERS_23_3_port
                           , S => n632, Z => n2447);
   U2958 : MUX2_X1 port map( A => REGISTERS_20_3_port, B => REGISTERS_22_3_port
                           , S => n632, Z => n2448);
   U2959 : MUX2_X1 port map( A => n2448, B => n2447, S => n665, Z => n2449);
   U2960 : MUX2_X1 port map( A => REGISTERS_17_3_port, B => REGISTERS_19_3_port
                           , S => n632, Z => n2450);
   U2961 : MUX2_X1 port map( A => REGISTERS_16_3_port, B => REGISTERS_18_3_port
                           , S => n632, Z => n2451);
   U2962 : MUX2_X1 port map( A => n2451, B => n2450, S => n665, Z => n2452);
   U2963 : MUX2_X1 port map( A => n2452, B => n2449, S => n592, Z => n2453);
   U2964 : MUX2_X1 port map( A => n2453, B => n2446, S => r3013_A_3_port, Z => 
                           n2454);
   U2965 : MUX2_X1 port map( A => REGISTERS_13_3_port, B => REGISTERS_15_3_port
                           , S => n631, Z => n2455);
   U2966 : MUX2_X1 port map( A => REGISTERS_12_3_port, B => REGISTERS_14_3_port
                           , S => n631, Z => n2456);
   U2967 : MUX2_X1 port map( A => n2456, B => n2455, S => n665, Z => n2457);
   U2968 : MUX2_X1 port map( A => REGISTERS_9_3_port, B => REGISTERS_11_3_port,
                           S => n631, Z => n2458);
   U2969 : MUX2_X1 port map( A => REGISTERS_8_3_port, B => REGISTERS_10_3_port,
                           S => n631, Z => n2459);
   U2970 : MUX2_X1 port map( A => n2459, B => n2458, S => n664, Z => n2460);
   U2971 : MUX2_X1 port map( A => n2460, B => n2457, S => n591, Z => n2461);
   U2972 : MUX2_X1 port map( A => REGISTERS_5_3_port, B => REGISTERS_7_3_port, 
                           S => n631, Z => n2462);
   U2973 : MUX2_X1 port map( A => REGISTERS_4_3_port, B => REGISTERS_6_3_port, 
                           S => n631, Z => n2463);
   U2974 : MUX2_X1 port map( A => n2463, B => n2462, S => n664, Z => n2464);
   U2975 : MUX2_X1 port map( A => REGISTERS_1_3_port, B => REGISTERS_3_3_port, 
                           S => n631, Z => n2465);
   U2976 : MUX2_X1 port map( A => REGISTERS_0_3_port, B => REGISTERS_2_3_port, 
                           S => n631, Z => n2466);
   U2977 : MUX2_X1 port map( A => n2466, B => n2465, S => n664, Z => n2467);
   U2978 : MUX2_X1 port map( A => n2467, B => n2464, S => n591, Z => n2468);
   U2979 : MUX2_X1 port map( A => n2468, B => n2461, S => r3013_A_3_port, Z => 
                           n2469);
   U2980 : MUX2_X1 port map( A => n2469, B => n2454, S => r3013_A_4_port, Z => 
                           n2470);
   U2981 : MUX2_X1 port map( A => n2470, B => n2439, S => ADD_RD2_5_port, Z => 
                           N4523);
   U2982 : MUX2_X1 port map( A => REGISTERS_37_4_port, B => REGISTERS_39_4_port
                           , S => n631, Z => n2471);
   U2983 : MUX2_X1 port map( A => REGISTERS_36_4_port, B => REGISTERS_38_4_port
                           , S => n631, Z => n2472);
   U2984 : MUX2_X1 port map( A => n2472, B => n2471, S => n664, Z => n2473);
   U2985 : MUX2_X1 port map( A => REGISTERS_33_4_port, B => REGISTERS_35_4_port
                           , S => n631, Z => n2474);
   U2986 : MUX2_X1 port map( A => REGISTERS_32_4_port, B => REGISTERS_34_4_port
                           , S => n631, Z => n2475);
   U2987 : MUX2_X1 port map( A => n2475, B => n2474, S => n664, Z => n2476);
   U2988 : MUX2_X1 port map( A => n2476, B => n2473, S => n591, Z => n2477);
   U2989 : MUX2_X1 port map( A => REGISTERS_29_4_port, B => REGISTERS_31_4_port
                           , S => n631, Z => n2478);
   U2990 : MUX2_X1 port map( A => REGISTERS_28_4_port, B => REGISTERS_30_4_port
                           , S => n631, Z => n2479);
   U2991 : MUX2_X1 port map( A => n2479, B => n2478, S => n664, Z => n2480);
   U2992 : MUX2_X1 port map( A => REGISTERS_25_4_port, B => REGISTERS_27_4_port
                           , S => n631, Z => n2481);
   U2993 : MUX2_X1 port map( A => REGISTERS_24_4_port, B => REGISTERS_26_4_port
                           , S => n630, Z => n2482);
   U2994 : MUX2_X1 port map( A => n2482, B => n2481, S => n664, Z => n2483);
   U2995 : MUX2_X1 port map( A => n2483, B => n2480, S => n591, Z => n2484);
   U2996 : MUX2_X1 port map( A => REGISTERS_21_4_port, B => REGISTERS_23_4_port
                           , S => n630, Z => n2485);
   U2997 : MUX2_X1 port map( A => REGISTERS_20_4_port, B => REGISTERS_22_4_port
                           , S => n630, Z => n2486);
   U2998 : MUX2_X1 port map( A => n2486, B => n2485, S => n664, Z => n2487);
   U2999 : MUX2_X1 port map( A => REGISTERS_17_4_port, B => REGISTERS_19_4_port
                           , S => n630, Z => n2488);
   U3000 : MUX2_X1 port map( A => REGISTERS_16_4_port, B => REGISTERS_18_4_port
                           , S => n630, Z => n2489);
   U3001 : MUX2_X1 port map( A => n2489, B => n2488, S => n664, Z => n2490);
   U3002 : MUX2_X1 port map( A => n2490, B => n2487, S => n591, Z => n2491);
   U3003 : MUX2_X1 port map( A => n2491, B => n2484, S => r3013_A_3_port, Z => 
                           n2492);
   U3004 : MUX2_X1 port map( A => REGISTERS_13_4_port, B => REGISTERS_15_4_port
                           , S => n630, Z => n2493);
   U3005 : MUX2_X1 port map( A => REGISTERS_12_4_port, B => REGISTERS_14_4_port
                           , S => n630, Z => n2494);
   U3006 : MUX2_X1 port map( A => n2494, B => n2493, S => n664, Z => n2495);
   U3007 : MUX2_X1 port map( A => REGISTERS_9_4_port, B => REGISTERS_11_4_port,
                           S => n630, Z => n2496);
   U3008 : MUX2_X1 port map( A => REGISTERS_8_4_port, B => REGISTERS_10_4_port,
                           S => n630, Z => n2497);
   U3009 : MUX2_X1 port map( A => n2497, B => n2496, S => n664, Z => n2498);
   U3010 : MUX2_X1 port map( A => n2498, B => n2495, S => n591, Z => n2499);
   U3011 : MUX2_X1 port map( A => REGISTERS_5_4_port, B => REGISTERS_7_4_port, 
                           S => n630, Z => n2500);
   U3012 : MUX2_X1 port map( A => REGISTERS_4_4_port, B => REGISTERS_6_4_port, 
                           S => n630, Z => n2501);
   U3013 : MUX2_X1 port map( A => n2501, B => n2500, S => n664, Z => n2502);
   U3014 : MUX2_X1 port map( A => REGISTERS_1_4_port, B => REGISTERS_3_4_port, 
                           S => n630, Z => n2503);
   U3015 : MUX2_X1 port map( A => REGISTERS_0_4_port, B => REGISTERS_2_4_port, 
                           S => n630, Z => n2504);
   U3016 : MUX2_X1 port map( A => n2504, B => n2503, S => n664, Z => n2505);
   U3017 : MUX2_X1 port map( A => n2505, B => n2502, S => n591, Z => n2506);
   U3018 : MUX2_X1 port map( A => n2506, B => n2499, S => r3013_A_3_port, Z => 
                           n2507);
   U3019 : MUX2_X1 port map( A => n2507, B => n2492, S => r3013_A_4_port, Z => 
                           n2508);
   U3020 : MUX2_X1 port map( A => n2508, B => n2477, S => ADD_RD2_5_port, Z => 
                           N4522);
   U3021 : MUX2_X1 port map( A => REGISTERS_37_5_port, B => REGISTERS_39_5_port
                           , S => n630, Z => n2509);
   U3022 : MUX2_X1 port map( A => REGISTERS_36_5_port, B => REGISTERS_38_5_port
                           , S => n630, Z => n2510);
   U3023 : MUX2_X1 port map( A => n2510, B => n2509, S => n664, Z => n2511);
   U3024 : MUX2_X1 port map( A => REGISTERS_33_5_port, B => REGISTERS_35_5_port
                           , S => n629, Z => n2512);
   U3025 : MUX2_X1 port map( A => REGISTERS_32_5_port, B => REGISTERS_34_5_port
                           , S => n629, Z => n2513);
   U3026 : MUX2_X1 port map( A => n2513, B => n2512, S => n664, Z => n2514);
   U3027 : MUX2_X1 port map( A => n2514, B => n2511, S => n591, Z => n2515);
   U3028 : MUX2_X1 port map( A => REGISTERS_29_5_port, B => REGISTERS_31_5_port
                           , S => n629, Z => n2516);
   U3029 : MUX2_X1 port map( A => REGISTERS_28_5_port, B => REGISTERS_30_5_port
                           , S => n629, Z => n2517);
   U3030 : MUX2_X1 port map( A => n2517, B => n2516, S => n663, Z => n2518);
   U3031 : MUX2_X1 port map( A => REGISTERS_25_5_port, B => REGISTERS_27_5_port
                           , S => n629, Z => n2519);
   U3032 : MUX2_X1 port map( A => REGISTERS_24_5_port, B => REGISTERS_26_5_port
                           , S => n629, Z => n2520);
   U3033 : MUX2_X1 port map( A => n2520, B => n2519, S => n663, Z => n2521);
   U3034 : MUX2_X1 port map( A => n2521, B => n2518, S => n591, Z => n2522);
   U3035 : MUX2_X1 port map( A => REGISTERS_21_5_port, B => REGISTERS_23_5_port
                           , S => n629, Z => n2523);
   U3036 : MUX2_X1 port map( A => REGISTERS_20_5_port, B => REGISTERS_22_5_port
                           , S => n629, Z => n2524);
   U3037 : MUX2_X1 port map( A => n2524, B => n2523, S => n663, Z => n2525);
   U3038 : MUX2_X1 port map( A => REGISTERS_17_5_port, B => REGISTERS_19_5_port
                           , S => n629, Z => n2526);
   U3039 : MUX2_X1 port map( A => REGISTERS_16_5_port, B => REGISTERS_18_5_port
                           , S => n629, Z => n2527);
   U3040 : MUX2_X1 port map( A => n2527, B => n2526, S => n663, Z => n2528);
   U3041 : MUX2_X1 port map( A => n2528, B => n2525, S => n591, Z => n2529);
   U3042 : MUX2_X1 port map( A => n2529, B => n2522, S => r3013_A_3_port, Z => 
                           n2530);
   U3043 : MUX2_X1 port map( A => REGISTERS_13_5_port, B => REGISTERS_15_5_port
                           , S => n629, Z => n2531);
   U3044 : MUX2_X1 port map( A => REGISTERS_12_5_port, B => REGISTERS_14_5_port
                           , S => n629, Z => n2532);
   U3045 : MUX2_X1 port map( A => n2532, B => n2531, S => n663, Z => n2533);
   U3046 : MUX2_X1 port map( A => REGISTERS_9_5_port, B => REGISTERS_11_5_port,
                           S => n629, Z => n2534);
   U3047 : MUX2_X1 port map( A => REGISTERS_8_5_port, B => REGISTERS_10_5_port,
                           S => n629, Z => n2535);
   U3048 : MUX2_X1 port map( A => n2535, B => n2534, S => n663, Z => n2536);
   U3049 : MUX2_X1 port map( A => n2536, B => n2533, S => n591, Z => n2537);
   U3050 : MUX2_X1 port map( A => REGISTERS_5_5_port, B => REGISTERS_7_5_port, 
                           S => n629, Z => n2538);
   U3051 : MUX2_X1 port map( A => REGISTERS_4_5_port, B => REGISTERS_6_5_port, 
                           S => n628, Z => n2539);
   U3052 : MUX2_X1 port map( A => n2539, B => n2538, S => n663, Z => n2540);
   U3053 : MUX2_X1 port map( A => REGISTERS_1_5_port, B => REGISTERS_3_5_port, 
                           S => n628, Z => n2541);
   U3054 : MUX2_X1 port map( A => REGISTERS_0_5_port, B => REGISTERS_2_5_port, 
                           S => n628, Z => n2542);
   U3055 : MUX2_X1 port map( A => n2542, B => n2541, S => n663, Z => n2543);
   U3056 : MUX2_X1 port map( A => n2543, B => n2540, S => n591, Z => n2544);
   U3057 : MUX2_X1 port map( A => n2544, B => n2537, S => r3013_A_3_port, Z => 
                           n2545);
   U3058 : MUX2_X1 port map( A => n2545, B => n2530, S => r3013_A_4_port, Z => 
                           n2546);
   U3059 : MUX2_X1 port map( A => n2546, B => n2515, S => ADD_RD2_5_port, Z => 
                           N4521);
   U3060 : MUX2_X1 port map( A => REGISTERS_37_6_port, B => REGISTERS_39_6_port
                           , S => n628, Z => n2547);
   U3061 : MUX2_X1 port map( A => REGISTERS_36_6_port, B => REGISTERS_38_6_port
                           , S => n628, Z => n2548);
   U3062 : MUX2_X1 port map( A => n2548, B => n2547, S => n663, Z => n2549);
   U3063 : MUX2_X1 port map( A => REGISTERS_33_6_port, B => REGISTERS_35_6_port
                           , S => n628, Z => n2550);
   U3064 : MUX2_X1 port map( A => REGISTERS_32_6_port, B => REGISTERS_34_6_port
                           , S => n628, Z => n2551);
   U3065 : MUX2_X1 port map( A => n2551, B => n2550, S => n663, Z => n2552);
   U3066 : MUX2_X1 port map( A => n2552, B => n2549, S => n591, Z => n2553);
   U3067 : MUX2_X1 port map( A => REGISTERS_29_6_port, B => REGISTERS_31_6_port
                           , S => n628, Z => n2554);
   U3068 : MUX2_X1 port map( A => REGISTERS_28_6_port, B => REGISTERS_30_6_port
                           , S => n628, Z => n2555);
   U3069 : MUX2_X1 port map( A => n2555, B => n2554, S => n663, Z => n2556);
   U3070 : MUX2_X1 port map( A => REGISTERS_25_6_port, B => REGISTERS_27_6_port
                           , S => n628, Z => n2557);
   U3071 : MUX2_X1 port map( A => REGISTERS_24_6_port, B => REGISTERS_26_6_port
                           , S => n628, Z => n2558);
   U3072 : MUX2_X1 port map( A => n2558, B => n2557, S => n663, Z => n2559);
   U3073 : MUX2_X1 port map( A => n2559, B => n2556, S => n590, Z => n2560);
   U3074 : MUX2_X1 port map( A => REGISTERS_21_6_port, B => REGISTERS_23_6_port
                           , S => n628, Z => n2561);
   U3075 : MUX2_X1 port map( A => REGISTERS_20_6_port, B => REGISTERS_22_6_port
                           , S => n628, Z => n2562);
   U3076 : MUX2_X1 port map( A => n2562, B => n2561, S => n663, Z => n2563);
   U3077 : MUX2_X1 port map( A => REGISTERS_17_6_port, B => REGISTERS_19_6_port
                           , S => n628, Z => n2564);
   U3078 : MUX2_X1 port map( A => REGISTERS_16_6_port, B => REGISTERS_18_6_port
                           , S => n628, Z => n2565);
   U3079 : MUX2_X1 port map( A => n2565, B => n2564, S => n663, Z => n2566);
   U3080 : MUX2_X1 port map( A => n2566, B => n2563, S => n590, Z => n2567);
   U3081 : MUX2_X1 port map( A => n2567, B => n2560, S => r3013_A_3_port, Z => 
                           n2568);
   U3082 : MUX2_X1 port map( A => REGISTERS_13_6_port, B => REGISTERS_15_6_port
                           , S => n627, Z => n2569);
   U3083 : MUX2_X1 port map( A => REGISTERS_12_6_port, B => REGISTERS_14_6_port
                           , S => n627, Z => n2570);
   U3084 : MUX2_X1 port map( A => n2570, B => n2569, S => n663, Z => n2571);
   U3085 : MUX2_X1 port map( A => REGISTERS_9_6_port, B => REGISTERS_11_6_port,
                           S => n627, Z => n2572);
   U3086 : MUX2_X1 port map( A => REGISTERS_8_6_port, B => REGISTERS_10_6_port,
                           S => n627, Z => n2573);
   U3087 : MUX2_X1 port map( A => n2573, B => n2572, S => n662, Z => n2574);
   U3088 : MUX2_X1 port map( A => n2574, B => n2571, S => n590, Z => n2575);
   U3089 : MUX2_X1 port map( A => REGISTERS_5_6_port, B => REGISTERS_7_6_port, 
                           S => n627, Z => n2576);
   U3090 : MUX2_X1 port map( A => REGISTERS_4_6_port, B => REGISTERS_6_6_port, 
                           S => n627, Z => n2577);
   U3091 : MUX2_X1 port map( A => n2577, B => n2576, S => n662, Z => n2578);
   U3092 : MUX2_X1 port map( A => REGISTERS_1_6_port, B => REGISTERS_3_6_port, 
                           S => n627, Z => n2579);
   U3093 : MUX2_X1 port map( A => REGISTERS_0_6_port, B => REGISTERS_2_6_port, 
                           S => n627, Z => n2580);
   U3094 : MUX2_X1 port map( A => n2580, B => n2579, S => n662, Z => n2581);
   U3095 : MUX2_X1 port map( A => n2581, B => n2578, S => n590, Z => n2582);
   U3096 : MUX2_X1 port map( A => n2582, B => n2575, S => r3013_A_3_port, Z => 
                           n2583);
   U3097 : MUX2_X1 port map( A => n2583, B => n2568, S => r3013_A_4_port, Z => 
                           n2584);
   U3098 : MUX2_X1 port map( A => n2584, B => n2553, S => ADD_RD2_5_port, Z => 
                           N4520);
   U3099 : MUX2_X1 port map( A => REGISTERS_37_7_port, B => REGISTERS_39_7_port
                           , S => n627, Z => n2585);
   U3100 : MUX2_X1 port map( A => REGISTERS_36_7_port, B => REGISTERS_38_7_port
                           , S => n627, Z => n2586);
   U3101 : MUX2_X1 port map( A => n2586, B => n2585, S => n662, Z => n2587);
   U3102 : MUX2_X1 port map( A => REGISTERS_33_7_port, B => REGISTERS_35_7_port
                           , S => n627, Z => n2588);
   U3103 : MUX2_X1 port map( A => REGISTERS_32_7_port, B => REGISTERS_34_7_port
                           , S => n627, Z => n2589);
   U3104 : MUX2_X1 port map( A => n2589, B => n2588, S => n662, Z => n2590);
   U3105 : MUX2_X1 port map( A => n2590, B => n2587, S => n590, Z => n2591);
   U3106 : MUX2_X1 port map( A => REGISTERS_29_7_port, B => REGISTERS_31_7_port
                           , S => n627, Z => n2592);
   U3107 : MUX2_X1 port map( A => REGISTERS_28_7_port, B => REGISTERS_30_7_port
                           , S => n627, Z => n2593);
   U3108 : MUX2_X1 port map( A => n2593, B => n2592, S => n662, Z => n2594);
   U3109 : MUX2_X1 port map( A => REGISTERS_25_7_port, B => REGISTERS_27_7_port
                           , S => n627, Z => n2595);
   U3110 : MUX2_X1 port map( A => REGISTERS_24_7_port, B => REGISTERS_26_7_port
                           , S => n626, Z => n2596);
   U3111 : MUX2_X1 port map( A => n2596, B => n2595, S => n662, Z => n2597);
   U3112 : MUX2_X1 port map( A => n2597, B => n2594, S => n590, Z => n2598);
   U3113 : MUX2_X1 port map( A => REGISTERS_21_7_port, B => REGISTERS_23_7_port
                           , S => n626, Z => n2599);
   U3114 : MUX2_X1 port map( A => REGISTERS_20_7_port, B => REGISTERS_22_7_port
                           , S => n626, Z => n2600);
   U3115 : MUX2_X1 port map( A => n2600, B => n2599, S => n662, Z => n2601);
   U3116 : MUX2_X1 port map( A => REGISTERS_17_7_port, B => REGISTERS_19_7_port
                           , S => n626, Z => n2602);
   U3117 : MUX2_X1 port map( A => REGISTERS_16_7_port, B => REGISTERS_18_7_port
                           , S => n626, Z => n2603);
   U3118 : MUX2_X1 port map( A => n2603, B => n2602, S => n662, Z => n2604);
   U3119 : MUX2_X1 port map( A => n2604, B => n2601, S => n590, Z => n2605);
   U3120 : MUX2_X1 port map( A => n2605, B => n2598, S => r3013_A_3_port, Z => 
                           n2606);
   U3121 : MUX2_X1 port map( A => REGISTERS_13_7_port, B => REGISTERS_15_7_port
                           , S => n626, Z => n2607);
   U3122 : MUX2_X1 port map( A => REGISTERS_12_7_port, B => REGISTERS_14_7_port
                           , S => n626, Z => n2608);
   U3123 : MUX2_X1 port map( A => n2608, B => n2607, S => n662, Z => n2609);
   U3124 : MUX2_X1 port map( A => REGISTERS_9_7_port, B => REGISTERS_11_7_port,
                           S => n626, Z => n2610);
   U3125 : MUX2_X1 port map( A => REGISTERS_8_7_port, B => REGISTERS_10_7_port,
                           S => n626, Z => n2611);
   U3126 : MUX2_X1 port map( A => n2611, B => n2610, S => n662, Z => n2612);
   U3127 : MUX2_X1 port map( A => n2612, B => n2609, S => n590, Z => n2613);
   U3128 : MUX2_X1 port map( A => REGISTERS_5_7_port, B => REGISTERS_7_7_port, 
                           S => n626, Z => n2614);
   U3129 : MUX2_X1 port map( A => REGISTERS_4_7_port, B => REGISTERS_6_7_port, 
                           S => n626, Z => n2615);
   U3130 : MUX2_X1 port map( A => n2615, B => n2614, S => n662, Z => n2616);
   U3131 : MUX2_X1 port map( A => REGISTERS_1_7_port, B => REGISTERS_3_7_port, 
                           S => n626, Z => n2617);
   U3132 : MUX2_X1 port map( A => REGISTERS_0_7_port, B => REGISTERS_2_7_port, 
                           S => n626, Z => n2618);
   U3133 : MUX2_X1 port map( A => n2618, B => n2617, S => n662, Z => n2619);
   U3134 : MUX2_X1 port map( A => n2619, B => n2616, S => n590, Z => n2620);
   U3135 : MUX2_X1 port map( A => n2620, B => n2613, S => r3013_A_3_port, Z => 
                           n2621);
   U3136 : MUX2_X1 port map( A => n2621, B => n2606, S => r3013_A_4_port, Z => 
                           n2622);
   U3137 : MUX2_X1 port map( A => n2622, B => n2591, S => ADD_RD2_5_port, Z => 
                           N4519);
   U3138 : MUX2_X1 port map( A => REGISTERS_37_8_port, B => REGISTERS_39_8_port
                           , S => n626, Z => n2623);
   U3139 : MUX2_X1 port map( A => REGISTERS_36_8_port, B => REGISTERS_38_8_port
                           , S => n626, Z => n2624);
   U3140 : MUX2_X1 port map( A => n2624, B => n2623, S => n662, Z => n2625);
   U3141 : MUX2_X1 port map( A => REGISTERS_33_8_port, B => REGISTERS_35_8_port
                           , S => n625, Z => n2626);
   U3142 : MUX2_X1 port map( A => REGISTERS_32_8_port, B => REGISTERS_34_8_port
                           , S => n625, Z => n2627);
   U3143 : MUX2_X1 port map( A => n2627, B => n2626, S => n662, Z => n2628);
   U3144 : MUX2_X1 port map( A => n2628, B => n2625, S => n590, Z => n2629);
   U3145 : MUX2_X1 port map( A => REGISTERS_29_8_port, B => REGISTERS_31_8_port
                           , S => n625, Z => n2630);
   U3146 : MUX2_X1 port map( A => REGISTERS_28_8_port, B => REGISTERS_30_8_port
                           , S => n625, Z => n2631);
   U3147 : MUX2_X1 port map( A => n2631, B => n2630, S => n661, Z => n2632);
   U3148 : MUX2_X1 port map( A => REGISTERS_25_8_port, B => REGISTERS_27_8_port
                           , S => n625, Z => n2633);
   U3149 : MUX2_X1 port map( A => REGISTERS_24_8_port, B => REGISTERS_26_8_port
                           , S => n625, Z => n2634);
   U3150 : MUX2_X1 port map( A => n2634, B => n2633, S => n661, Z => n2635);
   U3151 : MUX2_X1 port map( A => n2635, B => n2632, S => n590, Z => n2636);
   U3152 : MUX2_X1 port map( A => REGISTERS_21_8_port, B => REGISTERS_23_8_port
                           , S => n625, Z => n2637);
   U3153 : MUX2_X1 port map( A => REGISTERS_20_8_port, B => REGISTERS_22_8_port
                           , S => n625, Z => n2638);
   U3154 : MUX2_X1 port map( A => n2638, B => n2637, S => n661, Z => n2639);
   U3155 : MUX2_X1 port map( A => REGISTERS_17_8_port, B => REGISTERS_19_8_port
                           , S => n625, Z => n2640);
   U3156 : MUX2_X1 port map( A => REGISTERS_16_8_port, B => REGISTERS_18_8_port
                           , S => n625, Z => n2641);
   U3157 : MUX2_X1 port map( A => n2641, B => n2640, S => n661, Z => n2642);
   U3158 : MUX2_X1 port map( A => n2642, B => n2639, S => n590, Z => n2643);
   U3159 : MUX2_X1 port map( A => n2643, B => n2636, S => r3013_A_3_port, Z => 
                           n2644);
   U3160 : MUX2_X1 port map( A => REGISTERS_13_8_port, B => REGISTERS_15_8_port
                           , S => n625, Z => n2645);
   U3161 : MUX2_X1 port map( A => REGISTERS_12_8_port, B => REGISTERS_14_8_port
                           , S => n625, Z => n2646);
   U3162 : MUX2_X1 port map( A => n2646, B => n2645, S => n661, Z => n2647);
   U3163 : MUX2_X1 port map( A => REGISTERS_9_8_port, B => REGISTERS_11_8_port,
                           S => n625, Z => n2648);
   U3164 : MUX2_X1 port map( A => REGISTERS_8_8_port, B => REGISTERS_10_8_port,
                           S => n625, Z => n2649);
   U3165 : MUX2_X1 port map( A => n2649, B => n2648, S => n661, Z => n2650);
   U3166 : MUX2_X1 port map( A => n2650, B => n2647, S => n590, Z => n2651);
   U3167 : MUX2_X1 port map( A => REGISTERS_5_8_port, B => REGISTERS_7_8_port, 
                           S => n625, Z => n2652);
   U3168 : MUX2_X1 port map( A => REGISTERS_4_8_port, B => REGISTERS_6_8_port, 
                           S => n624, Z => n2653);
   U3169 : MUX2_X1 port map( A => n2653, B => n2652, S => n661, Z => n2654);
   U3170 : MUX2_X1 port map( A => REGISTERS_1_8_port, B => REGISTERS_3_8_port, 
                           S => n624, Z => n2655);
   U3171 : MUX2_X1 port map( A => REGISTERS_0_8_port, B => REGISTERS_2_8_port, 
                           S => n624, Z => n2656);
   U3172 : MUX2_X1 port map( A => n2656, B => n2655, S => n661, Z => n2657);
   U3173 : MUX2_X1 port map( A => n2657, B => n2654, S => n589, Z => n2658);
   U3174 : MUX2_X1 port map( A => n2658, B => n2651, S => r3013_A_3_port, Z => 
                           n2659);
   U3175 : MUX2_X1 port map( A => n2659, B => n2644, S => r3013_A_4_port, Z => 
                           n2660);
   U3176 : MUX2_X1 port map( A => n2660, B => n2629, S => ADD_RD2_5_port, Z => 
                           N4518);
   U3177 : MUX2_X1 port map( A => REGISTERS_37_9_port, B => REGISTERS_39_9_port
                           , S => n624, Z => n2661);
   U3178 : MUX2_X1 port map( A => REGISTERS_36_9_port, B => REGISTERS_38_9_port
                           , S => n624, Z => n2662);
   U3179 : MUX2_X1 port map( A => n2662, B => n2661, S => n661, Z => n2663);
   U3180 : MUX2_X1 port map( A => REGISTERS_33_9_port, B => REGISTERS_35_9_port
                           , S => n624, Z => n2664);
   U3181 : MUX2_X1 port map( A => REGISTERS_32_9_port, B => REGISTERS_34_9_port
                           , S => n624, Z => n2665);
   U3182 : MUX2_X1 port map( A => n2665, B => n2664, S => n661, Z => n2666);
   U3183 : MUX2_X1 port map( A => n2666, B => n2663, S => n589, Z => n2667);
   U3184 : MUX2_X1 port map( A => REGISTERS_29_9_port, B => REGISTERS_31_9_port
                           , S => n624, Z => n2668);
   U3185 : MUX2_X1 port map( A => REGISTERS_28_9_port, B => REGISTERS_30_9_port
                           , S => n624, Z => n2669);
   U3186 : MUX2_X1 port map( A => n2669, B => n2668, S => n661, Z => n2670);
   U3187 : MUX2_X1 port map( A => REGISTERS_25_9_port, B => REGISTERS_27_9_port
                           , S => n624, Z => n2671);
   U3188 : MUX2_X1 port map( A => REGISTERS_24_9_port, B => REGISTERS_26_9_port
                           , S => n624, Z => n2672);
   U3189 : MUX2_X1 port map( A => n2672, B => n2671, S => n661, Z => n2673);
   U3190 : MUX2_X1 port map( A => n2673, B => n2670, S => n589, Z => n2674);
   U3191 : MUX2_X1 port map( A => REGISTERS_21_9_port, B => REGISTERS_23_9_port
                           , S => n624, Z => n2675);
   U3192 : MUX2_X1 port map( A => REGISTERS_20_9_port, B => REGISTERS_22_9_port
                           , S => n624, Z => n2676);
   U3193 : MUX2_X1 port map( A => n2676, B => n2675, S => n661, Z => n2677);
   U3194 : MUX2_X1 port map( A => REGISTERS_17_9_port, B => REGISTERS_19_9_port
                           , S => n624, Z => n2678);
   U3195 : MUX2_X1 port map( A => REGISTERS_16_9_port, B => REGISTERS_18_9_port
                           , S => n624, Z => n2679);
   U3196 : MUX2_X1 port map( A => n2679, B => n2678, S => n661, Z => n2680);
   U3197 : MUX2_X1 port map( A => n2680, B => n2677, S => n589, Z => n2681);
   U3198 : MUX2_X1 port map( A => n2681, B => n2674, S => r3013_A_3_port, Z => 
                           n2682);
   U3199 : MUX2_X1 port map( A => REGISTERS_13_9_port, B => REGISTERS_15_9_port
                           , S => n623, Z => n2683);
   U3200 : MUX2_X1 port map( A => REGISTERS_12_9_port, B => REGISTERS_14_9_port
                           , S => n623, Z => n2684);
   U3201 : MUX2_X1 port map( A => n2684, B => n2683, S => n661, Z => n2685);
   U3202 : MUX2_X1 port map( A => REGISTERS_9_9_port, B => REGISTERS_11_9_port,
                           S => n623, Z => n2686);
   U3203 : MUX2_X1 port map( A => REGISTERS_8_9_port, B => REGISTERS_10_9_port,
                           S => n623, Z => n2687);
   U3204 : MUX2_X1 port map( A => n2687, B => n2686, S => n660, Z => n2688);
   U3205 : MUX2_X1 port map( A => n2688, B => n2685, S => n589, Z => n2689);
   U3206 : MUX2_X1 port map( A => REGISTERS_5_9_port, B => REGISTERS_7_9_port, 
                           S => n623, Z => n2690);
   U3207 : MUX2_X1 port map( A => REGISTERS_4_9_port, B => REGISTERS_6_9_port, 
                           S => n623, Z => n2691);
   U3208 : MUX2_X1 port map( A => n2691, B => n2690, S => n660, Z => n2692);
   U3209 : MUX2_X1 port map( A => REGISTERS_1_9_port, B => REGISTERS_3_9_port, 
                           S => n623, Z => n2693);
   U3210 : MUX2_X1 port map( A => REGISTERS_0_9_port, B => REGISTERS_2_9_port, 
                           S => n623, Z => n2694);
   U3211 : MUX2_X1 port map( A => n2694, B => n2693, S => n660, Z => n2695);
   U3212 : MUX2_X1 port map( A => n2695, B => n2692, S => n589, Z => n2696);
   U3213 : MUX2_X1 port map( A => n2696, B => n2689, S => r3013_A_3_port, Z => 
                           n2697);
   U3214 : MUX2_X1 port map( A => n2697, B => n2682, S => r3013_A_4_port, Z => 
                           n2698);
   U3215 : MUX2_X1 port map( A => n2698, B => n2667, S => ADD_RD2_5_port, Z => 
                           N4517);
   U3216 : MUX2_X1 port map( A => REGISTERS_37_10_port, B => 
                           REGISTERS_39_10_port, S => n623, Z => n2699);
   U3217 : MUX2_X1 port map( A => REGISTERS_36_10_port, B => 
                           REGISTERS_38_10_port, S => n623, Z => n2700);
   U3218 : MUX2_X1 port map( A => n2700, B => n2699, S => n660, Z => n2701);
   U3219 : MUX2_X1 port map( A => REGISTERS_33_10_port, B => 
                           REGISTERS_35_10_port, S => n623, Z => n2702);
   U3220 : MUX2_X1 port map( A => REGISTERS_32_10_port, B => 
                           REGISTERS_34_10_port, S => n623, Z => n2703);
   U3221 : MUX2_X1 port map( A => n2703, B => n2702, S => n660, Z => n2704);
   U3222 : MUX2_X1 port map( A => n2704, B => n2701, S => n589, Z => n2705);
   U3223 : MUX2_X1 port map( A => REGISTERS_29_10_port, B => 
                           REGISTERS_31_10_port, S => n623, Z => n2706);
   U3224 : MUX2_X1 port map( A => REGISTERS_28_10_port, B => 
                           REGISTERS_30_10_port, S => n623, Z => n2707);
   U3225 : MUX2_X1 port map( A => n2707, B => n2706, S => n660, Z => n2708);
   U3226 : MUX2_X1 port map( A => REGISTERS_25_10_port, B => 
                           REGISTERS_27_10_port, S => n623, Z => n2709);
   U3227 : MUX2_X1 port map( A => REGISTERS_24_10_port, B => 
                           REGISTERS_26_10_port, S => n622, Z => n2710);
   U3228 : MUX2_X1 port map( A => n2710, B => n2709, S => n660, Z => n2711);
   U3229 : MUX2_X1 port map( A => n2711, B => n2708, S => n589, Z => n2712);
   U3230 : MUX2_X1 port map( A => REGISTERS_21_10_port, B => 
                           REGISTERS_23_10_port, S => n622, Z => n2713);
   U3231 : MUX2_X1 port map( A => REGISTERS_20_10_port, B => 
                           REGISTERS_22_10_port, S => n622, Z => n2714);
   U3232 : MUX2_X1 port map( A => n2714, B => n2713, S => n660, Z => n2715);
   U3233 : MUX2_X1 port map( A => REGISTERS_17_10_port, B => 
                           REGISTERS_19_10_port, S => n622, Z => n2716);
   U3234 : MUX2_X1 port map( A => REGISTERS_16_10_port, B => 
                           REGISTERS_18_10_port, S => n622, Z => n2717);
   U3235 : MUX2_X1 port map( A => n2717, B => n2716, S => n660, Z => n2718);
   U3236 : MUX2_X1 port map( A => n2718, B => n2715, S => n589, Z => n2719);
   U3237 : MUX2_X1 port map( A => n2719, B => n2712, S => r3013_A_3_port, Z => 
                           n2720);
   U3238 : MUX2_X1 port map( A => REGISTERS_13_10_port, B => 
                           REGISTERS_15_10_port, S => n622, Z => n2721);
   U3239 : MUX2_X1 port map( A => REGISTERS_12_10_port, B => 
                           REGISTERS_14_10_port, S => n622, Z => n2722);
   U3240 : MUX2_X1 port map( A => n2722, B => n2721, S => n660, Z => n2723);
   U3241 : MUX2_X1 port map( A => REGISTERS_9_10_port, B => 
                           REGISTERS_11_10_port, S => n622, Z => n2724);
   U3242 : MUX2_X1 port map( A => REGISTERS_8_10_port, B => 
                           REGISTERS_10_10_port, S => n622, Z => n2725);
   U3243 : MUX2_X1 port map( A => n2725, B => n2724, S => n660, Z => n2726);
   U3244 : MUX2_X1 port map( A => n2726, B => n2723, S => n589, Z => n2727);
   U3245 : MUX2_X1 port map( A => REGISTERS_5_10_port, B => REGISTERS_7_10_port
                           , S => n622, Z => n2728);
   U3246 : MUX2_X1 port map( A => REGISTERS_4_10_port, B => REGISTERS_6_10_port
                           , S => n622, Z => n2729);
   U3247 : MUX2_X1 port map( A => n2729, B => n2728, S => n660, Z => n2730);
   U3248 : MUX2_X1 port map( A => REGISTERS_1_10_port, B => REGISTERS_3_10_port
                           , S => n622, Z => n2731);
   U3249 : MUX2_X1 port map( A => REGISTERS_0_10_port, B => REGISTERS_2_10_port
                           , S => n622, Z => n2732);
   U3250 : MUX2_X1 port map( A => n2732, B => n2731, S => n660, Z => n2733);
   U3251 : MUX2_X1 port map( A => n2733, B => n2730, S => n589, Z => n2734);
   U3252 : MUX2_X1 port map( A => n2734, B => n2727, S => r3013_A_3_port, Z => 
                           n2735);
   U3253 : MUX2_X1 port map( A => n2735, B => n2720, S => r3013_A_4_port, Z => 
                           n2736);
   U3254 : MUX2_X1 port map( A => n2736, B => n2705, S => ADD_RD2_5_port, Z => 
                           N4516);
   U3255 : MUX2_X1 port map( A => REGISTERS_37_11_port, B => 
                           REGISTERS_39_11_port, S => n622, Z => n2737);
   U3256 : MUX2_X1 port map( A => REGISTERS_36_11_port, B => 
                           REGISTERS_38_11_port, S => n622, Z => n2738);
   U3257 : MUX2_X1 port map( A => n2738, B => n2737, S => n660, Z => n2739);
   U3258 : MUX2_X1 port map( A => REGISTERS_33_11_port, B => 
                           REGISTERS_35_11_port, S => n621, Z => n2740);
   U3259 : MUX2_X1 port map( A => REGISTERS_32_11_port, B => 
                           REGISTERS_34_11_port, S => n621, Z => n2741);
   U3260 : MUX2_X1 port map( A => n2741, B => n2740, S => n660, Z => n2742);
   U3261 : MUX2_X1 port map( A => n2742, B => n2739, S => n589, Z => n2743);
   U3262 : MUX2_X1 port map( A => REGISTERS_29_11_port, B => 
                           REGISTERS_31_11_port, S => n621, Z => n2744);
   U3263 : MUX2_X1 port map( A => REGISTERS_28_11_port, B => 
                           REGISTERS_30_11_port, S => n621, Z => n2745);
   U3264 : MUX2_X1 port map( A => n2745, B => n2744, S => n659, Z => n2746);
   U3265 : MUX2_X1 port map( A => REGISTERS_25_11_port, B => 
                           REGISTERS_27_11_port, S => n621, Z => n2747);
   U3266 : MUX2_X1 port map( A => REGISTERS_24_11_port, B => 
                           REGISTERS_26_11_port, S => n621, Z => n2748);
   U3267 : MUX2_X1 port map( A => n2748, B => n2747, S => n659, Z => n2749);
   U3268 : MUX2_X1 port map( A => n2749, B => n2746, S => n589, Z => n2750);
   U3269 : MUX2_X1 port map( A => REGISTERS_21_11_port, B => 
                           REGISTERS_23_11_port, S => n621, Z => n2751);
   U3270 : MUX2_X1 port map( A => REGISTERS_20_11_port, B => 
                           REGISTERS_22_11_port, S => n621, Z => n2752);
   U3271 : MUX2_X1 port map( A => n2752, B => n2751, S => n659, Z => n2753);
   U3272 : MUX2_X1 port map( A => REGISTERS_17_11_port, B => 
                           REGISTERS_19_11_port, S => n621, Z => n2754);
   U3273 : MUX2_X1 port map( A => REGISTERS_16_11_port, B => 
                           REGISTERS_18_11_port, S => n621, Z => n2755);
   U3274 : MUX2_X1 port map( A => n2755, B => n2754, S => n659, Z => n2756);
   U3275 : MUX2_X1 port map( A => n2756, B => n2753, S => n588, Z => n2757);
   U3276 : MUX2_X1 port map( A => n2757, B => n2750, S => r3013_A_3_port, Z => 
                           n2758);
   U3277 : MUX2_X1 port map( A => REGISTERS_13_11_port, B => 
                           REGISTERS_15_11_port, S => n621, Z => n2759);
   U3278 : MUX2_X1 port map( A => REGISTERS_12_11_port, B => 
                           REGISTERS_14_11_port, S => n621, Z => n2760);
   U3279 : MUX2_X1 port map( A => n2760, B => n2759, S => n659, Z => n2761);
   U3280 : MUX2_X1 port map( A => REGISTERS_9_11_port, B => 
                           REGISTERS_11_11_port, S => n621, Z => n2762);
   U3281 : MUX2_X1 port map( A => REGISTERS_8_11_port, B => 
                           REGISTERS_10_11_port, S => n621, Z => n2763);
   U3282 : MUX2_X1 port map( A => n2763, B => n2762, S => n659, Z => n2764);
   U3283 : MUX2_X1 port map( A => n2764, B => n2761, S => n588, Z => n2765);
   U3284 : MUX2_X1 port map( A => REGISTERS_5_11_port, B => REGISTERS_7_11_port
                           , S => n621, Z => n2766);
   U3285 : MUX2_X1 port map( A => REGISTERS_4_11_port, B => REGISTERS_6_11_port
                           , S => n620, Z => n2767);
   U3286 : MUX2_X1 port map( A => n2767, B => n2766, S => n659, Z => n2768);
   U3287 : MUX2_X1 port map( A => REGISTERS_1_11_port, B => REGISTERS_3_11_port
                           , S => n620, Z => n2769);
   U3288 : MUX2_X1 port map( A => REGISTERS_0_11_port, B => REGISTERS_2_11_port
                           , S => n620, Z => n2770);
   U3289 : MUX2_X1 port map( A => n2770, B => n2769, S => n659, Z => n2771);
   U3290 : MUX2_X1 port map( A => n2771, B => n2768, S => n588, Z => n2772);
   U3291 : MUX2_X1 port map( A => n2772, B => n2765, S => r3013_A_3_port, Z => 
                           n2773);
   U3292 : MUX2_X1 port map( A => n2773, B => n2758, S => r3013_A_4_port, Z => 
                           n2774);
   U3293 : MUX2_X1 port map( A => n2774, B => n2743, S => ADD_RD2_5_port, Z => 
                           N4515);
   U3294 : MUX2_X1 port map( A => REGISTERS_37_12_port, B => 
                           REGISTERS_39_12_port, S => n620, Z => n2775);
   U3295 : MUX2_X1 port map( A => REGISTERS_36_12_port, B => 
                           REGISTERS_38_12_port, S => n620, Z => n2776);
   U3296 : MUX2_X1 port map( A => n2776, B => n2775, S => n659, Z => n2777);
   U3297 : MUX2_X1 port map( A => REGISTERS_33_12_port, B => 
                           REGISTERS_35_12_port, S => n620, Z => n2778);
   U3298 : MUX2_X1 port map( A => REGISTERS_32_12_port, B => 
                           REGISTERS_34_12_port, S => n620, Z => n2779);
   U3299 : MUX2_X1 port map( A => n2779, B => n2778, S => n659, Z => n2780);
   U3300 : MUX2_X1 port map( A => n2780, B => n2777, S => n588, Z => n2781);
   U3301 : MUX2_X1 port map( A => REGISTERS_29_12_port, B => 
                           REGISTERS_31_12_port, S => n620, Z => n2782);
   U3302 : MUX2_X1 port map( A => REGISTERS_28_12_port, B => 
                           REGISTERS_30_12_port, S => n620, Z => n2783);
   U3303 : MUX2_X1 port map( A => n2783, B => n2782, S => n659, Z => n2784);
   U3304 : MUX2_X1 port map( A => REGISTERS_25_12_port, B => 
                           REGISTERS_27_12_port, S => n620, Z => n2785);
   U3305 : MUX2_X1 port map( A => REGISTERS_24_12_port, B => 
                           REGISTERS_26_12_port, S => n620, Z => n2786);
   U3306 : MUX2_X1 port map( A => n2786, B => n2785, S => n659, Z => n2787);
   U3307 : MUX2_X1 port map( A => n2787, B => n2784, S => n588, Z => n2788);
   U3308 : MUX2_X1 port map( A => REGISTERS_21_12_port, B => 
                           REGISTERS_23_12_port, S => n620, Z => n2789);
   U3309 : MUX2_X1 port map( A => REGISTERS_20_12_port, B => 
                           REGISTERS_22_12_port, S => n620, Z => n2790);
   U3310 : MUX2_X1 port map( A => n2790, B => n2789, S => n659, Z => n2791);
   U3311 : MUX2_X1 port map( A => REGISTERS_17_12_port, B => 
                           REGISTERS_19_12_port, S => n620, Z => n2792);
   U3312 : MUX2_X1 port map( A => REGISTERS_16_12_port, B => 
                           REGISTERS_18_12_port, S => n620, Z => n2793);
   U3313 : MUX2_X1 port map( A => n2793, B => n2792, S => n659, Z => n2794);
   U3314 : MUX2_X1 port map( A => n2794, B => n2791, S => n588, Z => n2795);
   U3315 : MUX2_X1 port map( A => n2795, B => n2788, S => r3013_A_3_port, Z => 
                           n2796);
   U3316 : MUX2_X1 port map( A => REGISTERS_13_12_port, B => 
                           REGISTERS_15_12_port, S => n619, Z => n2797);
   U3317 : MUX2_X1 port map( A => REGISTERS_12_12_port, B => 
                           REGISTERS_14_12_port, S => n619, Z => n2798);
   U3318 : MUX2_X1 port map( A => n2798, B => n2797, S => n659, Z => n2799);
   U3319 : MUX2_X1 port map( A => REGISTERS_9_12_port, B => 
                           REGISTERS_11_12_port, S => n619, Z => n2800);
   U3320 : MUX2_X1 port map( A => REGISTERS_8_12_port, B => 
                           REGISTERS_10_12_port, S => n619, Z => n2801);
   U3321 : MUX2_X1 port map( A => n2801, B => n2800, S => n658, Z => n2802);
   U3322 : MUX2_X1 port map( A => n2802, B => n2799, S => n588, Z => n2803);
   U3323 : MUX2_X1 port map( A => REGISTERS_5_12_port, B => REGISTERS_7_12_port
                           , S => n619, Z => n2804);
   U3324 : MUX2_X1 port map( A => REGISTERS_4_12_port, B => REGISTERS_6_12_port
                           , S => n619, Z => n2805);
   U3325 : MUX2_X1 port map( A => n2805, B => n2804, S => n658, Z => n2806);
   U3326 : MUX2_X1 port map( A => REGISTERS_1_12_port, B => REGISTERS_3_12_port
                           , S => n619, Z => n2807);
   U3327 : MUX2_X1 port map( A => REGISTERS_0_12_port, B => REGISTERS_2_12_port
                           , S => n619, Z => n2808);
   U3328 : MUX2_X1 port map( A => n2808, B => n2807, S => n658, Z => n2809);
   U3329 : MUX2_X1 port map( A => n2809, B => n2806, S => n588, Z => n2810);
   U3330 : MUX2_X1 port map( A => n2810, B => n2803, S => r3013_A_3_port, Z => 
                           n2811);
   U3331 : MUX2_X1 port map( A => n2811, B => n2796, S => r3013_A_4_port, Z => 
                           n2812);
   U3332 : MUX2_X1 port map( A => n2812, B => n2781, S => ADD_RD2_5_port, Z => 
                           N4514);
   U3333 : MUX2_X1 port map( A => REGISTERS_37_13_port, B => 
                           REGISTERS_39_13_port, S => n619, Z => n2813);
   U3334 : MUX2_X1 port map( A => REGISTERS_36_13_port, B => 
                           REGISTERS_38_13_port, S => n619, Z => n2814);
   U3335 : MUX2_X1 port map( A => n2814, B => n2813, S => n658, Z => n2815);
   U3336 : MUX2_X1 port map( A => REGISTERS_33_13_port, B => 
                           REGISTERS_35_13_port, S => n619, Z => n2816);
   U3337 : MUX2_X1 port map( A => REGISTERS_32_13_port, B => 
                           REGISTERS_34_13_port, S => n619, Z => n2817);
   U3338 : MUX2_X1 port map( A => n2817, B => n2816, S => n658, Z => n2818);
   U3339 : MUX2_X1 port map( A => n2818, B => n2815, S => n588, Z => n2819);
   U3340 : MUX2_X1 port map( A => REGISTERS_29_13_port, B => 
                           REGISTERS_31_13_port, S => n619, Z => n2820);
   U3341 : MUX2_X1 port map( A => REGISTERS_28_13_port, B => 
                           REGISTERS_30_13_port, S => n619, Z => n2821);
   U3342 : MUX2_X1 port map( A => n2821, B => n2820, S => n658, Z => n2822);
   U3343 : MUX2_X1 port map( A => REGISTERS_25_13_port, B => 
                           REGISTERS_27_13_port, S => n619, Z => n2823);
   U3344 : MUX2_X1 port map( A => REGISTERS_24_13_port, B => 
                           REGISTERS_26_13_port, S => n618, Z => n2824);
   U3345 : MUX2_X1 port map( A => n2824, B => n2823, S => n658, Z => n2825);
   U3346 : MUX2_X1 port map( A => n2825, B => n2822, S => n588, Z => n2826);
   U3347 : MUX2_X1 port map( A => REGISTERS_21_13_port, B => 
                           REGISTERS_23_13_port, S => n618, Z => n2827);
   U3348 : MUX2_X1 port map( A => REGISTERS_20_13_port, B => 
                           REGISTERS_22_13_port, S => n618, Z => n2828);
   U3349 : MUX2_X1 port map( A => n2828, B => n2827, S => n658, Z => n2829);
   U3350 : MUX2_X1 port map( A => REGISTERS_17_13_port, B => 
                           REGISTERS_19_13_port, S => n618, Z => n2830);
   U3351 : MUX2_X1 port map( A => REGISTERS_16_13_port, B => 
                           REGISTERS_18_13_port, S => n618, Z => n2831);
   U3352 : MUX2_X1 port map( A => n2831, B => n2830, S => n658, Z => n2832);
   U3353 : MUX2_X1 port map( A => n2832, B => n2829, S => n588, Z => n2833);
   U3354 : MUX2_X1 port map( A => n2833, B => n2826, S => r3013_A_3_port, Z => 
                           n2834);
   U3355 : MUX2_X1 port map( A => REGISTERS_13_13_port, B => 
                           REGISTERS_15_13_port, S => n618, Z => n2835);
   U3356 : MUX2_X1 port map( A => REGISTERS_12_13_port, B => 
                           REGISTERS_14_13_port, S => n618, Z => n2836);
   U3357 : MUX2_X1 port map( A => n2836, B => n2835, S => n658, Z => n2837);
   U3358 : MUX2_X1 port map( A => REGISTERS_9_13_port, B => 
                           REGISTERS_11_13_port, S => n618, Z => n2838);
   U3359 : MUX2_X1 port map( A => REGISTERS_8_13_port, B => 
                           REGISTERS_10_13_port, S => n618, Z => n2839);
   U3360 : MUX2_X1 port map( A => n2839, B => n2838, S => n658, Z => n2840);
   U3361 : MUX2_X1 port map( A => n2840, B => n2837, S => n588, Z => n2841);
   U3362 : MUX2_X1 port map( A => REGISTERS_5_13_port, B => REGISTERS_7_13_port
                           , S => n618, Z => n2842);
   U3363 : MUX2_X1 port map( A => REGISTERS_4_13_port, B => REGISTERS_6_13_port
                           , S => n618, Z => n2843);
   U3364 : MUX2_X1 port map( A => n2843, B => n2842, S => n658, Z => n2844);
   U3365 : MUX2_X1 port map( A => REGISTERS_1_13_port, B => REGISTERS_3_13_port
                           , S => n618, Z => n2845);
   U3366 : MUX2_X1 port map( A => REGISTERS_0_13_port, B => REGISTERS_2_13_port
                           , S => n618, Z => n2846);
   U3367 : MUX2_X1 port map( A => n2846, B => n2845, S => n658, Z => n2847);
   U3368 : MUX2_X1 port map( A => n2847, B => n2844, S => n588, Z => n2848);
   U3369 : MUX2_X1 port map( A => n2848, B => n2841, S => r3013_A_3_port, Z => 
                           n2849);
   U3370 : MUX2_X1 port map( A => n2849, B => n2834, S => r3013_A_4_port, Z => 
                           n2850);
   U3371 : MUX2_X1 port map( A => n2850, B => n2819, S => ADD_RD2_5_port, Z => 
                           N4513);
   U3372 : MUX2_X1 port map( A => REGISTERS_37_14_port, B => 
                           REGISTERS_39_14_port, S => n618, Z => n2851);
   U3373 : MUX2_X1 port map( A => REGISTERS_36_14_port, B => 
                           REGISTERS_38_14_port, S => n618, Z => n2852);
   U3374 : MUX2_X1 port map( A => n2852, B => n2851, S => n658, Z => n2853);
   U3375 : MUX2_X1 port map( A => REGISTERS_33_14_port, B => 
                           REGISTERS_35_14_port, S => n617, Z => n2854);
   U3376 : MUX2_X1 port map( A => REGISTERS_32_14_port, B => 
                           REGISTERS_34_14_port, S => n617, Z => n2855);
   U3377 : MUX2_X1 port map( A => n2855, B => n2854, S => n658, Z => n2856);
   U3378 : MUX2_X1 port map( A => n2856, B => n2853, S => n587, Z => n2857);
   U3379 : MUX2_X1 port map( A => REGISTERS_29_14_port, B => 
                           REGISTERS_31_14_port, S => n617, Z => n2858);
   U3380 : MUX2_X1 port map( A => REGISTERS_28_14_port, B => 
                           REGISTERS_30_14_port, S => n617, Z => n2859);
   U3381 : MUX2_X1 port map( A => n2859, B => n2858, S => n657, Z => n2860);
   U3382 : MUX2_X1 port map( A => REGISTERS_25_14_port, B => 
                           REGISTERS_27_14_port, S => n617, Z => n2861);
   U3383 : MUX2_X1 port map( A => REGISTERS_24_14_port, B => 
                           REGISTERS_26_14_port, S => n617, Z => n2862);
   U3384 : MUX2_X1 port map( A => n2862, B => n2861, S => n657, Z => n2863);
   U3385 : MUX2_X1 port map( A => n2863, B => n2860, S => n587, Z => n2864);
   U3386 : MUX2_X1 port map( A => REGISTERS_21_14_port, B => 
                           REGISTERS_23_14_port, S => n617, Z => n2865);
   U3387 : MUX2_X1 port map( A => REGISTERS_20_14_port, B => 
                           REGISTERS_22_14_port, S => n617, Z => n2866);
   U3388 : MUX2_X1 port map( A => n2866, B => n2865, S => n657, Z => n2867);
   U3389 : MUX2_X1 port map( A => REGISTERS_17_14_port, B => 
                           REGISTERS_19_14_port, S => n617, Z => n2868);
   U3390 : MUX2_X1 port map( A => REGISTERS_16_14_port, B => 
                           REGISTERS_18_14_port, S => n617, Z => n2869);
   U3391 : MUX2_X1 port map( A => n2869, B => n2868, S => n657, Z => n2870);
   U3392 : MUX2_X1 port map( A => n2870, B => n2867, S => n587, Z => n2871);
   U3393 : MUX2_X1 port map( A => n2871, B => n2864, S => r3013_A_3_port, Z => 
                           n2872);
   U3394 : MUX2_X1 port map( A => REGISTERS_13_14_port, B => 
                           REGISTERS_15_14_port, S => n617, Z => n2873);
   U3395 : MUX2_X1 port map( A => REGISTERS_12_14_port, B => 
                           REGISTERS_14_14_port, S => n617, Z => n2874);
   U3396 : MUX2_X1 port map( A => n2874, B => n2873, S => n657, Z => n2875);
   U3397 : MUX2_X1 port map( A => REGISTERS_9_14_port, B => 
                           REGISTERS_11_14_port, S => n617, Z => n2876);
   U3398 : MUX2_X1 port map( A => REGISTERS_8_14_port, B => 
                           REGISTERS_10_14_port, S => n617, Z => n2877);
   U3399 : MUX2_X1 port map( A => n2877, B => n2876, S => n657, Z => n2878);
   U3400 : MUX2_X1 port map( A => n2878, B => n2875, S => n587, Z => n2879);
   U3401 : MUX2_X1 port map( A => REGISTERS_5_14_port, B => REGISTERS_7_14_port
                           , S => n617, Z => n2880);
   U3402 : MUX2_X1 port map( A => REGISTERS_4_14_port, B => REGISTERS_6_14_port
                           , S => n616, Z => n2881);
   U3403 : MUX2_X1 port map( A => n2881, B => n2880, S => n657, Z => n2882);
   U3404 : MUX2_X1 port map( A => REGISTERS_1_14_port, B => REGISTERS_3_14_port
                           , S => n616, Z => n2883);
   U3405 : MUX2_X1 port map( A => REGISTERS_0_14_port, B => REGISTERS_2_14_port
                           , S => n616, Z => n2884);
   U3406 : MUX2_X1 port map( A => n2884, B => n2883, S => n657, Z => n2885);
   U3407 : MUX2_X1 port map( A => n2885, B => n2882, S => n587, Z => n2886);
   U3408 : MUX2_X1 port map( A => n2886, B => n2879, S => r3013_A_3_port, Z => 
                           n2887);
   U3409 : MUX2_X1 port map( A => n2887, B => n2872, S => r3013_A_4_port, Z => 
                           n2888);
   U3410 : MUX2_X1 port map( A => n2888, B => n2857, S => ADD_RD2_5_port, Z => 
                           N4512);
   U3411 : MUX2_X1 port map( A => REGISTERS_37_15_port, B => 
                           REGISTERS_39_15_port, S => n616, Z => n2889);
   U3412 : MUX2_X1 port map( A => REGISTERS_36_15_port, B => 
                           REGISTERS_38_15_port, S => n616, Z => n2890);
   U3413 : MUX2_X1 port map( A => n2890, B => n2889, S => n657, Z => n2891);
   U3414 : MUX2_X1 port map( A => REGISTERS_33_15_port, B => 
                           REGISTERS_35_15_port, S => n616, Z => n2892);
   U3415 : MUX2_X1 port map( A => REGISTERS_32_15_port, B => 
                           REGISTERS_34_15_port, S => n616, Z => n2893);
   U3416 : MUX2_X1 port map( A => n2893, B => n2892, S => n657, Z => n2894);
   U3417 : MUX2_X1 port map( A => n2894, B => n2891, S => n587, Z => n2895);
   U3418 : MUX2_X1 port map( A => REGISTERS_29_15_port, B => 
                           REGISTERS_31_15_port, S => n616, Z => n2896);
   U3419 : MUX2_X1 port map( A => REGISTERS_28_15_port, B => 
                           REGISTERS_30_15_port, S => n616, Z => n2897);
   U3420 : MUX2_X1 port map( A => n2897, B => n2896, S => n657, Z => n2898);
   U3421 : MUX2_X1 port map( A => REGISTERS_25_15_port, B => 
                           REGISTERS_27_15_port, S => n616, Z => n2899);
   U3422 : MUX2_X1 port map( A => REGISTERS_24_15_port, B => 
                           REGISTERS_26_15_port, S => n616, Z => n2900);
   U3423 : MUX2_X1 port map( A => n2900, B => n2899, S => n657, Z => n2901);
   U3424 : MUX2_X1 port map( A => n2901, B => n2898, S => n587, Z => n2902);
   U3425 : MUX2_X1 port map( A => REGISTERS_21_15_port, B => 
                           REGISTERS_23_15_port, S => n616, Z => n2903);
   U3426 : MUX2_X1 port map( A => REGISTERS_20_15_port, B => 
                           REGISTERS_22_15_port, S => n616, Z => n2904);
   U3427 : MUX2_X1 port map( A => n2904, B => n2903, S => n657, Z => n2905);
   U3428 : MUX2_X1 port map( A => REGISTERS_17_15_port, B => 
                           REGISTERS_19_15_port, S => n616, Z => n2906);
   U3429 : MUX2_X1 port map( A => REGISTERS_16_15_port, B => 
                           REGISTERS_18_15_port, S => n616, Z => n2907);
   U3430 : MUX2_X1 port map( A => n2907, B => n2906, S => n657, Z => n2908);
   U3431 : MUX2_X1 port map( A => n2908, B => n2905, S => n587, Z => n2909);
   U3432 : MUX2_X1 port map( A => n2909, B => n2902, S => r3013_A_3_port, Z => 
                           n2910);
   U3433 : MUX2_X1 port map( A => REGISTERS_13_15_port, B => 
                           REGISTERS_15_15_port, S => n615, Z => n2911);
   U3434 : MUX2_X1 port map( A => REGISTERS_12_15_port, B => 
                           REGISTERS_14_15_port, S => n615, Z => n2912);
   U3435 : MUX2_X1 port map( A => n2912, B => n2911, S => n657, Z => n2913);
   U3436 : MUX2_X1 port map( A => REGISTERS_9_15_port, B => 
                           REGISTERS_11_15_port, S => n615, Z => n2914);
   U3437 : MUX2_X1 port map( A => REGISTERS_8_15_port, B => 
                           REGISTERS_10_15_port, S => n615, Z => n2915);
   U3438 : MUX2_X1 port map( A => n2915, B => n2914, S => n656, Z => n2916);
   U3439 : MUX2_X1 port map( A => n2916, B => n2913, S => n587, Z => n2917);
   U3440 : MUX2_X1 port map( A => REGISTERS_5_15_port, B => REGISTERS_7_15_port
                           , S => n615, Z => n2918);
   U3441 : MUX2_X1 port map( A => REGISTERS_4_15_port, B => REGISTERS_6_15_port
                           , S => n615, Z => n2919);
   U3442 : MUX2_X1 port map( A => n2919, B => n2918, S => n656, Z => n2920);
   U3443 : MUX2_X1 port map( A => REGISTERS_1_15_port, B => REGISTERS_3_15_port
                           , S => n615, Z => n2921);
   U3444 : MUX2_X1 port map( A => REGISTERS_0_15_port, B => REGISTERS_2_15_port
                           , S => n615, Z => n2922);
   U3445 : MUX2_X1 port map( A => n2922, B => n2921, S => n656, Z => n2923);
   U3446 : MUX2_X1 port map( A => n2923, B => n2920, S => n587, Z => n2924);
   U3447 : MUX2_X1 port map( A => n2924, B => n2917, S => r3013_A_3_port, Z => 
                           n2925);
   U3448 : MUX2_X1 port map( A => n2925, B => n2910, S => r3013_A_4_port, Z => 
                           n2926);
   U3449 : MUX2_X1 port map( A => n2926, B => n2895, S => ADD_RD2_5_port, Z => 
                           N4511);
   U3450 : MUX2_X1 port map( A => REGISTERS_37_16_port, B => 
                           REGISTERS_39_16_port, S => n615, Z => n2927);
   U3451 : MUX2_X1 port map( A => REGISTERS_36_16_port, B => 
                           REGISTERS_38_16_port, S => n615, Z => n2928);
   U3452 : MUX2_X1 port map( A => n2928, B => n2927, S => n656, Z => n2929);
   U3453 : MUX2_X1 port map( A => REGISTERS_33_16_port, B => 
                           REGISTERS_35_16_port, S => n615, Z => n2930);
   U3454 : MUX2_X1 port map( A => REGISTERS_32_16_port, B => 
                           REGISTERS_34_16_port, S => n615, Z => n2931);
   U3455 : MUX2_X1 port map( A => n2931, B => n2930, S => n656, Z => n2932);
   U3456 : MUX2_X1 port map( A => n2932, B => n2929, S => n587, Z => n2933);
   U3457 : MUX2_X1 port map( A => REGISTERS_29_16_port, B => 
                           REGISTERS_31_16_port, S => n615, Z => n2934);
   U3458 : MUX2_X1 port map( A => REGISTERS_28_16_port, B => 
                           REGISTERS_30_16_port, S => n615, Z => n2935);
   U3459 : MUX2_X1 port map( A => n2935, B => n2934, S => n656, Z => n2936);
   U3460 : MUX2_X1 port map( A => REGISTERS_25_16_port, B => 
                           REGISTERS_27_16_port, S => n615, Z => n2937);
   U3461 : MUX2_X1 port map( A => REGISTERS_24_16_port, B => 
                           REGISTERS_26_16_port, S => n614, Z => n2938);
   U3462 : MUX2_X1 port map( A => n2938, B => n2937, S => n656, Z => n2939);
   U3463 : MUX2_X1 port map( A => n2939, B => n2936, S => n587, Z => n2940);
   U3464 : MUX2_X1 port map( A => REGISTERS_21_16_port, B => 
                           REGISTERS_23_16_port, S => n614, Z => n2941);
   U3465 : MUX2_X1 port map( A => REGISTERS_20_16_port, B => 
                           REGISTERS_22_16_port, S => n614, Z => n2942);
   U3466 : MUX2_X1 port map( A => n2942, B => n2941, S => n656, Z => n2943);
   U3467 : MUX2_X1 port map( A => REGISTERS_17_16_port, B => 
                           REGISTERS_19_16_port, S => n614, Z => n2944);
   U3468 : MUX2_X1 port map( A => REGISTERS_16_16_port, B => 
                           REGISTERS_18_16_port, S => n614, Z => n2945);
   U3469 : MUX2_X1 port map( A => n2945, B => n2944, S => n656, Z => n2946);
   U3470 : MUX2_X1 port map( A => n2946, B => n2943, S => n587, Z => n2947);
   U3471 : MUX2_X1 port map( A => n2947, B => n2940, S => r3013_A_3_port, Z => 
                           n2948);
   U3472 : MUX2_X1 port map( A => REGISTERS_13_16_port, B => 
                           REGISTERS_15_16_port, S => n614, Z => n2949);
   U3473 : MUX2_X1 port map( A => REGISTERS_12_16_port, B => 
                           REGISTERS_14_16_port, S => n614, Z => n2950);
   U3474 : MUX2_X1 port map( A => n2950, B => n2949, S => n656, Z => n2951);
   U3475 : MUX2_X1 port map( A => REGISTERS_9_16_port, B => 
                           REGISTERS_11_16_port, S => n614, Z => n2952);
   U3476 : MUX2_X1 port map( A => REGISTERS_8_16_port, B => 
                           REGISTERS_10_16_port, S => n614, Z => n2953);
   U3477 : MUX2_X1 port map( A => n2953, B => n2952, S => n656, Z => n2954);
   U3478 : MUX2_X1 port map( A => n2954, B => n2951, S => n586, Z => n2955);
   U3479 : MUX2_X1 port map( A => REGISTERS_5_16_port, B => REGISTERS_7_16_port
                           , S => n614, Z => n2956);
   U3480 : MUX2_X1 port map( A => REGISTERS_4_16_port, B => REGISTERS_6_16_port
                           , S => n614, Z => n2957);
   U3481 : MUX2_X1 port map( A => n2957, B => n2956, S => n656, Z => n2958);
   U3482 : MUX2_X1 port map( A => REGISTERS_1_16_port, B => REGISTERS_3_16_port
                           , S => n614, Z => n2959);
   U3483 : MUX2_X1 port map( A => REGISTERS_0_16_port, B => REGISTERS_2_16_port
                           , S => n614, Z => n2960);
   U3484 : MUX2_X1 port map( A => n2960, B => n2959, S => n656, Z => n2961);
   U3485 : MUX2_X1 port map( A => n2961, B => n2958, S => n586, Z => n2962);
   U3486 : MUX2_X1 port map( A => n2962, B => n2955, S => r3013_A_3_port, Z => 
                           n2963);
   U3487 : MUX2_X1 port map( A => n2963, B => n2948, S => r3013_A_4_port, Z => 
                           n2964);
   U3488 : MUX2_X1 port map( A => n2964, B => n2933, S => ADD_RD2_5_port, Z => 
                           N4510);
   U3489 : MUX2_X1 port map( A => REGISTERS_37_17_port, B => 
                           REGISTERS_39_17_port, S => n614, Z => n2965);
   U3490 : MUX2_X1 port map( A => REGISTERS_36_17_port, B => 
                           REGISTERS_38_17_port, S => n614, Z => n2966);
   U3491 : MUX2_X1 port map( A => n2966, B => n2965, S => n656, Z => n2967);
   U3492 : MUX2_X1 port map( A => REGISTERS_33_17_port, B => 
                           REGISTERS_35_17_port, S => n613, Z => n2968);
   U3493 : MUX2_X1 port map( A => REGISTERS_32_17_port, B => 
                           REGISTERS_34_17_port, S => n613, Z => n2969);
   U3494 : MUX2_X1 port map( A => n2969, B => n2968, S => n656, Z => n2970);
   U3495 : MUX2_X1 port map( A => n2970, B => n2967, S => n586, Z => n2971);
   U3496 : MUX2_X1 port map( A => REGISTERS_29_17_port, B => 
                           REGISTERS_31_17_port, S => n613, Z => n2972);
   U3497 : MUX2_X1 port map( A => REGISTERS_28_17_port, B => 
                           REGISTERS_30_17_port, S => n613, Z => n2973);
   U3498 : MUX2_X1 port map( A => n2973, B => n2972, S => n655, Z => n2974);
   U3499 : MUX2_X1 port map( A => REGISTERS_25_17_port, B => 
                           REGISTERS_27_17_port, S => n613, Z => n2975);
   U3500 : MUX2_X1 port map( A => REGISTERS_24_17_port, B => 
                           REGISTERS_26_17_port, S => n613, Z => n2976);
   U3501 : MUX2_X1 port map( A => n2976, B => n2975, S => n655, Z => n2977);
   U3502 : MUX2_X1 port map( A => n2977, B => n2974, S => n586, Z => n2978);
   U3503 : MUX2_X1 port map( A => REGISTERS_21_17_port, B => 
                           REGISTERS_23_17_port, S => n613, Z => n2979);
   U3504 : MUX2_X1 port map( A => REGISTERS_20_17_port, B => 
                           REGISTERS_22_17_port, S => n613, Z => n2980);
   U3505 : MUX2_X1 port map( A => n2980, B => n2979, S => n655, Z => n2981);
   U3506 : MUX2_X1 port map( A => REGISTERS_17_17_port, B => 
                           REGISTERS_19_17_port, S => n613, Z => n2982);
   U3507 : MUX2_X1 port map( A => REGISTERS_16_17_port, B => 
                           REGISTERS_18_17_port, S => n613, Z => n2983);
   U3508 : MUX2_X1 port map( A => n2983, B => n2982, S => n655, Z => n2984);
   U3509 : MUX2_X1 port map( A => n2984, B => n2981, S => n586, Z => n2985);
   U3510 : MUX2_X1 port map( A => n2985, B => n2978, S => r3013_A_3_port, Z => 
                           n2986);
   U3511 : MUX2_X1 port map( A => REGISTERS_13_17_port, B => 
                           REGISTERS_15_17_port, S => n613, Z => n2987);
   U3512 : MUX2_X1 port map( A => REGISTERS_12_17_port, B => 
                           REGISTERS_14_17_port, S => n613, Z => n2988);
   U3513 : MUX2_X1 port map( A => n2988, B => n2987, S => n655, Z => n2989);
   U3514 : MUX2_X1 port map( A => REGISTERS_9_17_port, B => 
                           REGISTERS_11_17_port, S => n613, Z => n2990);
   U3515 : MUX2_X1 port map( A => REGISTERS_8_17_port, B => 
                           REGISTERS_10_17_port, S => n613, Z => n2991);
   U3516 : MUX2_X1 port map( A => n2991, B => n2990, S => n655, Z => n2992);
   U3517 : MUX2_X1 port map( A => n2992, B => n2989, S => n586, Z => n2993);
   U3518 : MUX2_X1 port map( A => REGISTERS_5_17_port, B => REGISTERS_7_17_port
                           , S => n613, Z => n2994);
   U3519 : MUX2_X1 port map( A => REGISTERS_4_17_port, B => REGISTERS_6_17_port
                           , S => n612, Z => n2995);
   U3520 : MUX2_X1 port map( A => n2995, B => n2994, S => n655, Z => n2996);
   U3521 : MUX2_X1 port map( A => REGISTERS_1_17_port, B => REGISTERS_3_17_port
                           , S => n612, Z => n2997);
   U3522 : MUX2_X1 port map( A => REGISTERS_0_17_port, B => REGISTERS_2_17_port
                           , S => n612, Z => n2998);
   U3523 : MUX2_X1 port map( A => n2998, B => n2997, S => n655, Z => n2999);
   U3524 : MUX2_X1 port map( A => n2999, B => n2996, S => n586, Z => n3000);
   U3525 : MUX2_X1 port map( A => n3000, B => n2993, S => r3013_A_3_port, Z => 
                           n3001);
   U3526 : MUX2_X1 port map( A => n3001, B => n2986, S => r3013_A_4_port, Z => 
                           n3002);
   U3527 : MUX2_X1 port map( A => n3002, B => n2971, S => ADD_RD2_5_port, Z => 
                           N4509);
   U3528 : MUX2_X1 port map( A => REGISTERS_37_18_port, B => 
                           REGISTERS_39_18_port, S => n612, Z => n3003);
   U3529 : MUX2_X1 port map( A => REGISTERS_36_18_port, B => 
                           REGISTERS_38_18_port, S => n612, Z => n3004);
   U3530 : MUX2_X1 port map( A => n3004, B => n3003, S => n655, Z => n3005);
   U3531 : MUX2_X1 port map( A => REGISTERS_33_18_port, B => 
                           REGISTERS_35_18_port, S => n612, Z => n3006);
   U3532 : MUX2_X1 port map( A => REGISTERS_32_18_port, B => 
                           REGISTERS_34_18_port, S => n612, Z => n3007);
   U3533 : MUX2_X1 port map( A => n3007, B => n3006, S => n655, Z => n3008);
   U3534 : MUX2_X1 port map( A => n3008, B => n3005, S => n586, Z => n3009);
   U3535 : MUX2_X1 port map( A => REGISTERS_29_18_port, B => 
                           REGISTERS_31_18_port, S => n612, Z => n3010);
   U3536 : MUX2_X1 port map( A => REGISTERS_28_18_port, B => 
                           REGISTERS_30_18_port, S => n612, Z => n3011);
   U3537 : MUX2_X1 port map( A => n3011, B => n3010, S => n655, Z => n3012);
   U3538 : MUX2_X1 port map( A => REGISTERS_25_18_port, B => 
                           REGISTERS_27_18_port, S => n612, Z => n3013);
   U3539 : MUX2_X1 port map( A => REGISTERS_24_18_port, B => 
                           REGISTERS_26_18_port, S => n612, Z => n3014);
   U3540 : MUX2_X1 port map( A => n3014, B => n3013, S => n655, Z => n3015);
   U3541 : MUX2_X1 port map( A => n3015, B => n3012, S => n586, Z => n3016);
   U3542 : MUX2_X1 port map( A => REGISTERS_21_18_port, B => 
                           REGISTERS_23_18_port, S => n612, Z => n3017);
   U3543 : MUX2_X1 port map( A => REGISTERS_20_18_port, B => 
                           REGISTERS_22_18_port, S => n612, Z => n3018);
   U3544 : MUX2_X1 port map( A => n3018, B => n3017, S => n655, Z => n3019);
   U3545 : MUX2_X1 port map( A => REGISTERS_17_18_port, B => 
                           REGISTERS_19_18_port, S => n612, Z => n3020);
   U3546 : MUX2_X1 port map( A => REGISTERS_16_18_port, B => 
                           REGISTERS_18_18_port, S => n612, Z => n3021);
   U3547 : MUX2_X1 port map( A => n3021, B => n3020, S => n655, Z => n3022);
   U3548 : MUX2_X1 port map( A => n3022, B => n3019, S => n586, Z => n3023);
   U3549 : MUX2_X1 port map( A => n3023, B => n3016, S => r3013_A_3_port, Z => 
                           n3024);
   U3550 : MUX2_X1 port map( A => REGISTERS_13_18_port, B => 
                           REGISTERS_15_18_port, S => n611, Z => n3025);
   U3551 : MUX2_X1 port map( A => REGISTERS_12_18_port, B => 
                           REGISTERS_14_18_port, S => n611, Z => n3026);
   U3552 : MUX2_X1 port map( A => n3026, B => n3025, S => n655, Z => n3027);
   U3553 : MUX2_X1 port map( A => REGISTERS_9_18_port, B => 
                           REGISTERS_11_18_port, S => n611, Z => n3028);
   U3554 : MUX2_X1 port map( A => REGISTERS_8_18_port, B => 
                           REGISTERS_10_18_port, S => n611, Z => n3029);
   U3555 : MUX2_X1 port map( A => n3029, B => n3028, S => n654, Z => n3030);
   U3556 : MUX2_X1 port map( A => n3030, B => n3027, S => n586, Z => n3031);
   U3557 : MUX2_X1 port map( A => REGISTERS_5_18_port, B => REGISTERS_7_18_port
                           , S => n611, Z => n3032);
   U3558 : MUX2_X1 port map( A => REGISTERS_4_18_port, B => REGISTERS_6_18_port
                           , S => n611, Z => n3033);
   U3559 : MUX2_X1 port map( A => n3033, B => n3032, S => n654, Z => n3034);
   U3560 : MUX2_X1 port map( A => REGISTERS_1_18_port, B => REGISTERS_3_18_port
                           , S => n611, Z => n3035);
   U3561 : MUX2_X1 port map( A => REGISTERS_0_18_port, B => REGISTERS_2_18_port
                           , S => n611, Z => n3036);
   U3562 : MUX2_X1 port map( A => n3036, B => n3035, S => n654, Z => n3037);
   U3563 : MUX2_X1 port map( A => n3037, B => n3034, S => n586, Z => n3038);
   U3564 : MUX2_X1 port map( A => n3038, B => n3031, S => r3013_A_3_port, Z => 
                           n3039);
   U3565 : MUX2_X1 port map( A => n3039, B => n3024, S => r3013_A_4_port, Z => 
                           n3040);
   U3566 : MUX2_X1 port map( A => n3040, B => n3009, S => ADD_RD2_5_port, Z => 
                           N4508);
   U3567 : MUX2_X1 port map( A => REGISTERS_37_19_port, B => 
                           REGISTERS_39_19_port, S => n611, Z => n3041);
   U3568 : MUX2_X1 port map( A => REGISTERS_36_19_port, B => 
                           REGISTERS_38_19_port, S => n611, Z => n3042);
   U3569 : MUX2_X1 port map( A => n3042, B => n3041, S => n654, Z => n3043);
   U3570 : MUX2_X1 port map( A => REGISTERS_33_19_port, B => 
                           REGISTERS_35_19_port, S => n611, Z => n3044);
   U3571 : MUX2_X1 port map( A => REGISTERS_32_19_port, B => 
                           REGISTERS_34_19_port, S => n611, Z => n3045);
   U3572 : MUX2_X1 port map( A => n3045, B => n3044, S => n654, Z => n3046);
   U3573 : MUX2_X1 port map( A => n3046, B => n3043, S => n586, Z => n3047);
   U3574 : MUX2_X1 port map( A => REGISTERS_29_19_port, B => 
                           REGISTERS_31_19_port, S => n611, Z => n3048);
   U3575 : MUX2_X1 port map( A => REGISTERS_28_19_port, B => 
                           REGISTERS_30_19_port, S => n611, Z => n3049);
   U3576 : MUX2_X1 port map( A => n3049, B => n3048, S => n654, Z => n3050);
   U3577 : MUX2_X1 port map( A => REGISTERS_25_19_port, B => 
                           REGISTERS_27_19_port, S => n611, Z => n3051);
   U3578 : MUX2_X1 port map( A => REGISTERS_24_19_port, B => 
                           REGISTERS_26_19_port, S => n610, Z => n3052);
   U3579 : MUX2_X1 port map( A => n3052, B => n3051, S => n654, Z => n3053);
   U3580 : MUX2_X1 port map( A => n3053, B => n3050, S => n585, Z => n3054);
   U3581 : MUX2_X1 port map( A => REGISTERS_21_19_port, B => 
                           REGISTERS_23_19_port, S => n610, Z => n3055);
   U3582 : MUX2_X1 port map( A => REGISTERS_20_19_port, B => 
                           REGISTERS_22_19_port, S => n610, Z => n3056);
   U3583 : MUX2_X1 port map( A => n3056, B => n3055, S => n654, Z => n3057);
   U3584 : MUX2_X1 port map( A => REGISTERS_17_19_port, B => 
                           REGISTERS_19_19_port, S => n610, Z => n3058);
   U3585 : MUX2_X1 port map( A => REGISTERS_16_19_port, B => 
                           REGISTERS_18_19_port, S => n610, Z => n3059);
   U3586 : MUX2_X1 port map( A => n3059, B => n3058, S => n654, Z => n3060);
   U3587 : MUX2_X1 port map( A => n3060, B => n3057, S => n585, Z => n3061);
   U3588 : MUX2_X1 port map( A => n3061, B => n3054, S => r3013_A_3_port, Z => 
                           n3062);
   U3589 : MUX2_X1 port map( A => REGISTERS_13_19_port, B => 
                           REGISTERS_15_19_port, S => n610, Z => n3063);
   U3590 : MUX2_X1 port map( A => REGISTERS_12_19_port, B => 
                           REGISTERS_14_19_port, S => n610, Z => n3064);
   U3591 : MUX2_X1 port map( A => n3064, B => n3063, S => n654, Z => n3065);
   U3592 : MUX2_X1 port map( A => REGISTERS_9_19_port, B => 
                           REGISTERS_11_19_port, S => n610, Z => n3066);
   U3593 : MUX2_X1 port map( A => REGISTERS_8_19_port, B => 
                           REGISTERS_10_19_port, S => n610, Z => n3067);
   U3594 : MUX2_X1 port map( A => n3067, B => n3066, S => n654, Z => n3068);
   U3595 : MUX2_X1 port map( A => n3068, B => n3065, S => n585, Z => n3069);
   U3596 : MUX2_X1 port map( A => REGISTERS_5_19_port, B => REGISTERS_7_19_port
                           , S => n610, Z => n3070);
   U3597 : MUX2_X1 port map( A => REGISTERS_4_19_port, B => REGISTERS_6_19_port
                           , S => n610, Z => n3071);
   U3598 : MUX2_X1 port map( A => n3071, B => n3070, S => n654, Z => n3072);
   U3599 : MUX2_X1 port map( A => REGISTERS_1_19_port, B => REGISTERS_3_19_port
                           , S => n610, Z => n3073);
   U3600 : MUX2_X1 port map( A => REGISTERS_0_19_port, B => REGISTERS_2_19_port
                           , S => n610, Z => n3074);
   U3601 : MUX2_X1 port map( A => n3074, B => n3073, S => n654, Z => n3075);
   U3602 : MUX2_X1 port map( A => n3075, B => n3072, S => n585, Z => n3076);
   U3603 : MUX2_X1 port map( A => n3076, B => n3069, S => r3013_A_3_port, Z => 
                           n3077);
   U3604 : MUX2_X1 port map( A => n3077, B => n3062, S => r3013_A_4_port, Z => 
                           n3078);
   U3605 : MUX2_X1 port map( A => n3078, B => n3047, S => ADD_RD2_5_port, Z => 
                           N4507);
   U3606 : MUX2_X1 port map( A => REGISTERS_37_20_port, B => 
                           REGISTERS_39_20_port, S => n610, Z => n3079);
   U3607 : MUX2_X1 port map( A => REGISTERS_36_20_port, B => 
                           REGISTERS_38_20_port, S => n610, Z => n3080);
   U3608 : MUX2_X1 port map( A => n3080, B => n3079, S => n654, Z => n3081);
   U3609 : MUX2_X1 port map( A => REGISTERS_33_20_port, B => 
                           REGISTERS_35_20_port, S => n609, Z => n3082);
   U3610 : MUX2_X1 port map( A => REGISTERS_32_20_port, B => 
                           REGISTERS_34_20_port, S => n609, Z => n3083);
   U3611 : MUX2_X1 port map( A => n3083, B => n3082, S => n654, Z => n3084);
   U3612 : MUX2_X1 port map( A => n3084, B => n3081, S => n585, Z => n3085);
   U3613 : MUX2_X1 port map( A => REGISTERS_29_20_port, B => 
                           REGISTERS_31_20_port, S => n609, Z => n3086);
   U3614 : MUX2_X1 port map( A => REGISTERS_28_20_port, B => 
                           REGISTERS_30_20_port, S => n609, Z => n3087);
   U3615 : MUX2_X1 port map( A => n3087, B => n3086, S => n653, Z => n3088);
   U3616 : MUX2_X1 port map( A => REGISTERS_25_20_port, B => 
                           REGISTERS_27_20_port, S => n609, Z => n3089);
   U3617 : MUX2_X1 port map( A => REGISTERS_24_20_port, B => 
                           REGISTERS_26_20_port, S => n609, Z => n3090);
   U3618 : MUX2_X1 port map( A => n3090, B => n3089, S => n653, Z => n3091);
   U3619 : MUX2_X1 port map( A => n3091, B => n3088, S => n585, Z => n3092);
   U3620 : MUX2_X1 port map( A => REGISTERS_21_20_port, B => 
                           REGISTERS_23_20_port, S => n609, Z => n3093);
   U3621 : MUX2_X1 port map( A => REGISTERS_20_20_port, B => 
                           REGISTERS_22_20_port, S => n609, Z => n3094);
   U3622 : MUX2_X1 port map( A => n3094, B => n3093, S => n653, Z => n3095);
   U3623 : MUX2_X1 port map( A => REGISTERS_17_20_port, B => 
                           REGISTERS_19_20_port, S => n609, Z => n3096);
   U3624 : MUX2_X1 port map( A => REGISTERS_16_20_port, B => 
                           REGISTERS_18_20_port, S => n609, Z => n3097);
   U3625 : MUX2_X1 port map( A => n3097, B => n3096, S => n653, Z => n3098);
   U3626 : MUX2_X1 port map( A => n3098, B => n3095, S => n585, Z => n3099);
   U3627 : MUX2_X1 port map( A => n3099, B => n3092, S => r3013_A_3_port, Z => 
                           n3100);
   U3628 : MUX2_X1 port map( A => REGISTERS_13_20_port, B => 
                           REGISTERS_15_20_port, S => n609, Z => n3101);
   U3629 : MUX2_X1 port map( A => REGISTERS_12_20_port, B => 
                           REGISTERS_14_20_port, S => n609, Z => n3102);
   U3630 : MUX2_X1 port map( A => n3102, B => n3101, S => n653, Z => n3103);
   U3631 : MUX2_X1 port map( A => REGISTERS_9_20_port, B => 
                           REGISTERS_11_20_port, S => n609, Z => n3104);
   U3632 : MUX2_X1 port map( A => REGISTERS_8_20_port, B => 
                           REGISTERS_10_20_port, S => n609, Z => n3105);
   U3633 : MUX2_X1 port map( A => n3105, B => n3104, S => n653, Z => n3106);
   U3634 : MUX2_X1 port map( A => n3106, B => n3103, S => n585, Z => n3107);
   U3635 : MUX2_X1 port map( A => REGISTERS_5_20_port, B => REGISTERS_7_20_port
                           , S => n609, Z => n3108);
   U3636 : MUX2_X1 port map( A => REGISTERS_4_20_port, B => REGISTERS_6_20_port
                           , S => n608, Z => n3109);
   U3637 : MUX2_X1 port map( A => n3109, B => n3108, S => n653, Z => n3110);
   U3638 : MUX2_X1 port map( A => REGISTERS_1_20_port, B => REGISTERS_3_20_port
                           , S => n608, Z => n3111);
   U3639 : MUX2_X1 port map( A => REGISTERS_0_20_port, B => REGISTERS_2_20_port
                           , S => n608, Z => n3112);
   U3640 : MUX2_X1 port map( A => n3112, B => n3111, S => n653, Z => n3113);
   U3641 : MUX2_X1 port map( A => n3113, B => n3110, S => n585, Z => n3114);
   U3642 : MUX2_X1 port map( A => n3114, B => n3107, S => r3013_A_3_port, Z => 
                           n3115);
   U3643 : MUX2_X1 port map( A => n3115, B => n3100, S => r3013_A_4_port, Z => 
                           n3116);
   U3644 : MUX2_X1 port map( A => n3116, B => n3085, S => ADD_RD2_5_port, Z => 
                           N4506);
   U3645 : MUX2_X1 port map( A => REGISTERS_37_21_port, B => 
                           REGISTERS_39_21_port, S => n608, Z => n3117);
   U3646 : MUX2_X1 port map( A => REGISTERS_36_21_port, B => 
                           REGISTERS_38_21_port, S => n608, Z => n3118);
   U3647 : MUX2_X1 port map( A => n3118, B => n3117, S => n653, Z => n3119);
   U3648 : MUX2_X1 port map( A => REGISTERS_33_21_port, B => 
                           REGISTERS_35_21_port, S => n608, Z => n3120);
   U3649 : MUX2_X1 port map( A => REGISTERS_32_21_port, B => 
                           REGISTERS_34_21_port, S => n608, Z => n3121);
   U3650 : MUX2_X1 port map( A => n3121, B => n3120, S => n653, Z => n3122);
   U3651 : MUX2_X1 port map( A => n3122, B => n3119, S => n585, Z => n3123);
   U3652 : MUX2_X1 port map( A => REGISTERS_29_21_port, B => 
                           REGISTERS_31_21_port, S => n608, Z => n3124);
   U3653 : MUX2_X1 port map( A => REGISTERS_28_21_port, B => 
                           REGISTERS_30_21_port, S => n608, Z => n3125);
   U3654 : MUX2_X1 port map( A => n3125, B => n3124, S => n653, Z => n3126);
   U3655 : MUX2_X1 port map( A => REGISTERS_25_21_port, B => 
                           REGISTERS_27_21_port, S => n608, Z => n3127);
   U3656 : MUX2_X1 port map( A => REGISTERS_24_21_port, B => 
                           REGISTERS_26_21_port, S => n608, Z => n3128);
   U3657 : MUX2_X1 port map( A => n3128, B => n3127, S => n653, Z => n3129);
   U3658 : MUX2_X1 port map( A => n3129, B => n3126, S => n585, Z => n3130);
   U3659 : MUX2_X1 port map( A => REGISTERS_21_21_port, B => 
                           REGISTERS_23_21_port, S => n608, Z => n3131);
   U3660 : MUX2_X1 port map( A => REGISTERS_20_21_port, B => 
                           REGISTERS_22_21_port, S => n608, Z => n3132);
   U3661 : MUX2_X1 port map( A => n3132, B => n3131, S => n653, Z => n3133);
   U3662 : MUX2_X1 port map( A => REGISTERS_17_21_port, B => 
                           REGISTERS_19_21_port, S => n608, Z => n3134);
   U3663 : MUX2_X1 port map( A => REGISTERS_16_21_port, B => 
                           REGISTERS_18_21_port, S => n608, Z => n3135);
   U3664 : MUX2_X1 port map( A => n3135, B => n3134, S => n653, Z => n3136);
   U3665 : MUX2_X1 port map( A => n3136, B => n3133, S => n585, Z => n3137);
   U3666 : MUX2_X1 port map( A => n3137, B => n3130, S => r3013_A_3_port, Z => 
                           n3138);
   U3667 : MUX2_X1 port map( A => REGISTERS_13_21_port, B => 
                           REGISTERS_15_21_port, S => n607, Z => n3139);
   U3668 : MUX2_X1 port map( A => REGISTERS_12_21_port, B => 
                           REGISTERS_14_21_port, S => n607, Z => n3140);
   U3669 : MUX2_X1 port map( A => n3140, B => n3139, S => n653, Z => n3141);
   U3670 : MUX2_X1 port map( A => REGISTERS_9_21_port, B => 
                           REGISTERS_11_21_port, S => n607, Z => n3142);
   U3671 : MUX2_X1 port map( A => REGISTERS_8_21_port, B => 
                           REGISTERS_10_21_port, S => n607, Z => n3143);
   U3672 : MUX2_X1 port map( A => n3143, B => n3142, S => n652, Z => n3144);
   U3673 : MUX2_X1 port map( A => n3144, B => n3141, S => n585, Z => n3145);
   U3674 : MUX2_X1 port map( A => REGISTERS_5_21_port, B => REGISTERS_7_21_port
                           , S => n607, Z => n3146);
   U3675 : MUX2_X1 port map( A => REGISTERS_4_21_port, B => REGISTERS_6_21_port
                           , S => n607, Z => n3147);
   U3676 : MUX2_X1 port map( A => n3147, B => n3146, S => n652, Z => n3148);
   U3677 : MUX2_X1 port map( A => REGISTERS_1_21_port, B => REGISTERS_3_21_port
                           , S => n607, Z => n3149);
   U3678 : MUX2_X1 port map( A => REGISTERS_0_21_port, B => REGISTERS_2_21_port
                           , S => n607, Z => n3150);
   U3679 : MUX2_X1 port map( A => n3150, B => n3149, S => n652, Z => n3151);
   U3680 : MUX2_X1 port map( A => n3151, B => n3148, S => n584, Z => n3152);
   U3681 : MUX2_X1 port map( A => n3152, B => n3145, S => r3013_A_3_port, Z => 
                           n3153);
   U3682 : MUX2_X1 port map( A => n3153, B => n3138, S => r3013_A_4_port, Z => 
                           n3154);
   U3683 : MUX2_X1 port map( A => n3154, B => n3123, S => ADD_RD2_5_port, Z => 
                           N4505);
   U3684 : MUX2_X1 port map( A => REGISTERS_37_22_port, B => 
                           REGISTERS_39_22_port, S => n607, Z => n3155);
   U3685 : MUX2_X1 port map( A => REGISTERS_36_22_port, B => 
                           REGISTERS_38_22_port, S => n607, Z => n3156);
   U3686 : MUX2_X1 port map( A => n3156, B => n3155, S => n652, Z => n3157);
   U3687 : MUX2_X1 port map( A => REGISTERS_33_22_port, B => 
                           REGISTERS_35_22_port, S => n607, Z => n3158);
   U3688 : MUX2_X1 port map( A => REGISTERS_32_22_port, B => 
                           REGISTERS_34_22_port, S => n607, Z => n3159);
   U3689 : MUX2_X1 port map( A => n3159, B => n3158, S => n652, Z => n3160);
   U3690 : MUX2_X1 port map( A => n3160, B => n3157, S => n584, Z => n3161);
   U3691 : MUX2_X1 port map( A => REGISTERS_29_22_port, B => 
                           REGISTERS_31_22_port, S => n607, Z => n3162);
   U3692 : MUX2_X1 port map( A => REGISTERS_28_22_port, B => 
                           REGISTERS_30_22_port, S => n607, Z => n3163);
   U3693 : MUX2_X1 port map( A => n3163, B => n3162, S => n652, Z => n3164);
   U3694 : MUX2_X1 port map( A => REGISTERS_25_22_port, B => 
                           REGISTERS_27_22_port, S => n607, Z => n3165);
   U3695 : MUX2_X1 port map( A => REGISTERS_24_22_port, B => 
                           REGISTERS_26_22_port, S => n606, Z => n3166);
   U3696 : MUX2_X1 port map( A => n3166, B => n3165, S => n652, Z => n3167);
   U3697 : MUX2_X1 port map( A => n3167, B => n3164, S => n584, Z => n3168);
   U3698 : MUX2_X1 port map( A => REGISTERS_21_22_port, B => 
                           REGISTERS_23_22_port, S => n606, Z => n3169);
   U3699 : MUX2_X1 port map( A => REGISTERS_20_22_port, B => 
                           REGISTERS_22_22_port, S => n606, Z => n3170);
   U3700 : MUX2_X1 port map( A => n3170, B => n3169, S => n652, Z => n3171);
   U3701 : MUX2_X1 port map( A => REGISTERS_17_22_port, B => 
                           REGISTERS_19_22_port, S => n606, Z => n3172);
   U3702 : MUX2_X1 port map( A => REGISTERS_16_22_port, B => 
                           REGISTERS_18_22_port, S => n606, Z => n3173);
   U3703 : MUX2_X1 port map( A => n3173, B => n3172, S => n652, Z => n3174);
   U3704 : MUX2_X1 port map( A => n3174, B => n3171, S => n584, Z => n3175);
   U3705 : MUX2_X1 port map( A => n3175, B => n3168, S => r3013_A_3_port, Z => 
                           n3176);
   U3706 : MUX2_X1 port map( A => REGISTERS_13_22_port, B => 
                           REGISTERS_15_22_port, S => n606, Z => n3177);
   U3707 : MUX2_X1 port map( A => REGISTERS_12_22_port, B => 
                           REGISTERS_14_22_port, S => n606, Z => n3178);
   U3708 : MUX2_X1 port map( A => n3178, B => n3177, S => n652, Z => n3179);
   U3709 : MUX2_X1 port map( A => REGISTERS_9_22_port, B => 
                           REGISTERS_11_22_port, S => n606, Z => n3180);
   U3710 : MUX2_X1 port map( A => REGISTERS_8_22_port, B => 
                           REGISTERS_10_22_port, S => n606, Z => n3181);
   U3711 : MUX2_X1 port map( A => n3181, B => n3180, S => n652, Z => n3182);
   U3712 : MUX2_X1 port map( A => n3182, B => n3179, S => n584, Z => n3183);
   U3713 : MUX2_X1 port map( A => REGISTERS_5_22_port, B => REGISTERS_7_22_port
                           , S => n606, Z => n3184);
   U3714 : MUX2_X1 port map( A => REGISTERS_4_22_port, B => REGISTERS_6_22_port
                           , S => n606, Z => n3185);
   U3715 : MUX2_X1 port map( A => n3185, B => n3184, S => n652, Z => n3186);
   U3716 : MUX2_X1 port map( A => REGISTERS_1_22_port, B => REGISTERS_3_22_port
                           , S => n606, Z => n3187);
   U3717 : MUX2_X1 port map( A => REGISTERS_0_22_port, B => REGISTERS_2_22_port
                           , S => n606, Z => n3188);
   U3718 : MUX2_X1 port map( A => n3188, B => n3187, S => n652, Z => n3189);
   U3719 : MUX2_X1 port map( A => n3189, B => n3186, S => n584, Z => n3190);
   U3720 : MUX2_X1 port map( A => n3190, B => n3183, S => r3013_A_3_port, Z => 
                           n3191);
   U3721 : MUX2_X1 port map( A => n3191, B => n3176, S => r3013_A_4_port, Z => 
                           n3192);
   U3722 : MUX2_X1 port map( A => n3192, B => n3161, S => ADD_RD2_5_port, Z => 
                           N4504);
   U3723 : MUX2_X1 port map( A => REGISTERS_37_23_port, B => 
                           REGISTERS_39_23_port, S => n606, Z => n3193);
   U3724 : MUX2_X1 port map( A => REGISTERS_36_23_port, B => 
                           REGISTERS_38_23_port, S => n606, Z => n3194);
   U3725 : MUX2_X1 port map( A => n3194, B => n3193, S => n652, Z => n3195);
   U3726 : MUX2_X1 port map( A => REGISTERS_33_23_port, B => 
                           REGISTERS_35_23_port, S => n605, Z => n3196);
   U3727 : MUX2_X1 port map( A => REGISTERS_32_23_port, B => 
                           REGISTERS_34_23_port, S => n605, Z => n3197);
   U3728 : MUX2_X1 port map( A => n3197, B => n3196, S => n652, Z => n3198);
   U3729 : MUX2_X1 port map( A => n3198, B => n3195, S => n584, Z => n3199);
   U3730 : MUX2_X1 port map( A => REGISTERS_29_23_port, B => 
                           REGISTERS_31_23_port, S => n605, Z => n3200);
   U3731 : MUX2_X1 port map( A => REGISTERS_28_23_port, B => 
                           REGISTERS_30_23_port, S => n605, Z => n3201);
   U3732 : MUX2_X1 port map( A => n3201, B => n3200, S => n651, Z => n3202);
   U3733 : MUX2_X1 port map( A => REGISTERS_25_23_port, B => 
                           REGISTERS_27_23_port, S => n605, Z => n3203);
   U3734 : MUX2_X1 port map( A => REGISTERS_24_23_port, B => 
                           REGISTERS_26_23_port, S => n605, Z => n3204);
   U3735 : MUX2_X1 port map( A => n3204, B => n3203, S => n651, Z => n3205);
   U3736 : MUX2_X1 port map( A => n3205, B => n3202, S => n584, Z => n3206);
   U3737 : MUX2_X1 port map( A => REGISTERS_21_23_port, B => 
                           REGISTERS_23_23_port, S => n605, Z => n3207);
   U3738 : MUX2_X1 port map( A => REGISTERS_20_23_port, B => 
                           REGISTERS_22_23_port, S => n605, Z => n3208);
   U3739 : MUX2_X1 port map( A => n3208, B => n3207, S => n651, Z => n3209);
   U3740 : MUX2_X1 port map( A => REGISTERS_17_23_port, B => 
                           REGISTERS_19_23_port, S => n605, Z => n3210);
   U3741 : MUX2_X1 port map( A => REGISTERS_16_23_port, B => 
                           REGISTERS_18_23_port, S => n605, Z => n3211);
   U3742 : MUX2_X1 port map( A => n3211, B => n3210, S => n651, Z => n3212);
   U3743 : MUX2_X1 port map( A => n3212, B => n3209, S => n584, Z => n3213);
   U3744 : MUX2_X1 port map( A => n3213, B => n3206, S => r3013_A_3_port, Z => 
                           n3214);
   U3745 : MUX2_X1 port map( A => REGISTERS_13_23_port, B => 
                           REGISTERS_15_23_port, S => n605, Z => n3215);
   U3746 : MUX2_X1 port map( A => REGISTERS_12_23_port, B => 
                           REGISTERS_14_23_port, S => n605, Z => n3216);
   U3747 : MUX2_X1 port map( A => n3216, B => n3215, S => n651, Z => n3217);
   U3748 : MUX2_X1 port map( A => REGISTERS_9_23_port, B => 
                           REGISTERS_11_23_port, S => n605, Z => n3218);
   U3749 : MUX2_X1 port map( A => REGISTERS_8_23_port, B => 
                           REGISTERS_10_23_port, S => n605, Z => n3219);
   U3750 : MUX2_X1 port map( A => n3219, B => n3218, S => n651, Z => n3220);
   U3751 : MUX2_X1 port map( A => n3220, B => n3217, S => n584, Z => n3221);
   U3752 : MUX2_X1 port map( A => REGISTERS_5_23_port, B => REGISTERS_7_23_port
                           , S => n605, Z => n3222);
   U3753 : MUX2_X1 port map( A => REGISTERS_4_23_port, B => REGISTERS_6_23_port
                           , S => n604, Z => n3223);
   U3754 : MUX2_X1 port map( A => n3223, B => n3222, S => n651, Z => n3224);
   U3755 : MUX2_X1 port map( A => REGISTERS_1_23_port, B => REGISTERS_3_23_port
                           , S => n604, Z => n3225);
   U3756 : MUX2_X1 port map( A => REGISTERS_0_23_port, B => REGISTERS_2_23_port
                           , S => n604, Z => n3226);
   U3757 : MUX2_X1 port map( A => n3226, B => n3225, S => n651, Z => n3227);
   U3758 : MUX2_X1 port map( A => n3227, B => n3224, S => n584, Z => n3228);
   U3759 : MUX2_X1 port map( A => n3228, B => n3221, S => r3013_A_3_port, Z => 
                           n3229);
   U3760 : MUX2_X1 port map( A => n3229, B => n3214, S => r3013_A_4_port, Z => 
                           n3230);
   U3761 : MUX2_X1 port map( A => n3230, B => n3199, S => ADD_RD2_5_port, Z => 
                           N4503);
   U3762 : MUX2_X1 port map( A => REGISTERS_37_24_port, B => 
                           REGISTERS_39_24_port, S => n604, Z => n3231);
   U3763 : MUX2_X1 port map( A => REGISTERS_36_24_port, B => 
                           REGISTERS_38_24_port, S => n604, Z => n3232);
   U3764 : MUX2_X1 port map( A => n3232, B => n3231, S => n651, Z => n3233);
   U3765 : MUX2_X1 port map( A => REGISTERS_33_24_port, B => 
                           REGISTERS_35_24_port, S => n604, Z => n3234);
   U3766 : MUX2_X1 port map( A => REGISTERS_32_24_port, B => 
                           REGISTERS_34_24_port, S => n604, Z => n3235);
   U3767 : MUX2_X1 port map( A => n3235, B => n3234, S => n651, Z => n3236);
   U3768 : MUX2_X1 port map( A => n3236, B => n3233, S => n584, Z => n3237);
   U3769 : MUX2_X1 port map( A => REGISTERS_29_24_port, B => 
                           REGISTERS_31_24_port, S => n604, Z => n3238);
   U3770 : MUX2_X1 port map( A => REGISTERS_28_24_port, B => 
                           REGISTERS_30_24_port, S => n604, Z => n3239);
   U3771 : MUX2_X1 port map( A => n3239, B => n3238, S => n651, Z => n3240);
   U3772 : MUX2_X1 port map( A => REGISTERS_25_24_port, B => 
                           REGISTERS_27_24_port, S => n604, Z => n3241);
   U3773 : MUX2_X1 port map( A => REGISTERS_24_24_port, B => 
                           REGISTERS_26_24_port, S => n604, Z => n3242);
   U3774 : MUX2_X1 port map( A => n3242, B => n3241, S => n651, Z => n3243);
   U3775 : MUX2_X1 port map( A => n3243, B => n3240, S => n584, Z => n3244);
   U3776 : MUX2_X1 port map( A => REGISTERS_21_24_port, B => 
                           REGISTERS_23_24_port, S => n604, Z => n3245);
   U3777 : MUX2_X1 port map( A => REGISTERS_20_24_port, B => 
                           REGISTERS_22_24_port, S => n604, Z => n3246);
   U3778 : MUX2_X1 port map( A => n3246, B => n3245, S => n651, Z => n3247);
   U3779 : MUX2_X1 port map( A => REGISTERS_17_24_port, B => 
                           REGISTERS_19_24_port, S => n604, Z => n3248);
   U3780 : MUX2_X1 port map( A => REGISTERS_16_24_port, B => 
                           REGISTERS_18_24_port, S => n604, Z => n3249);
   U3781 : MUX2_X1 port map( A => n3249, B => n3248, S => n651, Z => n3250);
   U3782 : MUX2_X1 port map( A => n3250, B => n3247, S => n583, Z => n3251);
   U3783 : MUX2_X1 port map( A => n3251, B => n3244, S => r3013_A_3_port, Z => 
                           n3252);
   U3784 : MUX2_X1 port map( A => REGISTERS_13_24_port, B => 
                           REGISTERS_15_24_port, S => n603, Z => n3253);
   U3785 : MUX2_X1 port map( A => REGISTERS_12_24_port, B => 
                           REGISTERS_14_24_port, S => n603, Z => n3254);
   U3786 : MUX2_X1 port map( A => n3254, B => n3253, S => n651, Z => n3255);
   U3787 : MUX2_X1 port map( A => REGISTERS_9_24_port, B => 
                           REGISTERS_11_24_port, S => n603, Z => n3256);
   U3788 : MUX2_X1 port map( A => REGISTERS_8_24_port, B => 
                           REGISTERS_10_24_port, S => n603, Z => n3257);
   U3789 : MUX2_X1 port map( A => n3257, B => n3256, S => n650, Z => n3258);
   U3790 : MUX2_X1 port map( A => n3258, B => n3255, S => n583, Z => n3259);
   U3791 : MUX2_X1 port map( A => REGISTERS_5_24_port, B => REGISTERS_7_24_port
                           , S => n603, Z => n3260);
   U3792 : MUX2_X1 port map( A => REGISTERS_4_24_port, B => REGISTERS_6_24_port
                           , S => n603, Z => n3261);
   U3793 : MUX2_X1 port map( A => n3261, B => n3260, S => n650, Z => n3262);
   U3794 : MUX2_X1 port map( A => REGISTERS_1_24_port, B => REGISTERS_3_24_port
                           , S => n603, Z => n3263);
   U3795 : MUX2_X1 port map( A => REGISTERS_0_24_port, B => REGISTERS_2_24_port
                           , S => n603, Z => n3264);
   U3796 : MUX2_X1 port map( A => n3264, B => n3263, S => n650, Z => n3265);
   U3797 : MUX2_X1 port map( A => n3265, B => n3262, S => n583, Z => n3266);
   U3798 : MUX2_X1 port map( A => n3266, B => n3259, S => r3013_A_3_port, Z => 
                           n3267);
   U3799 : MUX2_X1 port map( A => n3267, B => n3252, S => r3013_A_4_port, Z => 
                           n3268);
   U3800 : MUX2_X1 port map( A => n3268, B => n3237, S => ADD_RD2_5_port, Z => 
                           N4502);
   U3801 : MUX2_X1 port map( A => REGISTERS_37_25_port, B => 
                           REGISTERS_39_25_port, S => n603, Z => n3269);
   U3802 : MUX2_X1 port map( A => REGISTERS_36_25_port, B => 
                           REGISTERS_38_25_port, S => n603, Z => n3270);
   U3803 : MUX2_X1 port map( A => n3270, B => n3269, S => n650, Z => n3271);
   U3804 : MUX2_X1 port map( A => REGISTERS_33_25_port, B => 
                           REGISTERS_35_25_port, S => n603, Z => n3272);
   U3805 : MUX2_X1 port map( A => REGISTERS_32_25_port, B => 
                           REGISTERS_34_25_port, S => n603, Z => n3273);
   U3806 : MUX2_X1 port map( A => n3273, B => n3272, S => n650, Z => n3274);
   U3807 : MUX2_X1 port map( A => n3274, B => n3271, S => n583, Z => n3275);
   U3808 : MUX2_X1 port map( A => REGISTERS_29_25_port, B => 
                           REGISTERS_31_25_port, S => n603, Z => n3276);
   U3809 : MUX2_X1 port map( A => REGISTERS_28_25_port, B => 
                           REGISTERS_30_25_port, S => n603, Z => n3277);
   U3810 : MUX2_X1 port map( A => n3277, B => n3276, S => n650, Z => n3278);
   U3811 : MUX2_X1 port map( A => REGISTERS_25_25_port, B => 
                           REGISTERS_27_25_port, S => n603, Z => n3279);
   U3812 : MUX2_X1 port map( A => REGISTERS_24_25_port, B => 
                           REGISTERS_26_25_port, S => n602, Z => n3280);
   U3813 : MUX2_X1 port map( A => n3280, B => n3279, S => n650, Z => n3281);
   U3814 : MUX2_X1 port map( A => n3281, B => n3278, S => n583, Z => n3282);
   U3815 : MUX2_X1 port map( A => REGISTERS_21_25_port, B => 
                           REGISTERS_23_25_port, S => n602, Z => n3283);
   U3816 : MUX2_X1 port map( A => REGISTERS_20_25_port, B => 
                           REGISTERS_22_25_port, S => n602, Z => n3284);
   U3817 : MUX2_X1 port map( A => n3284, B => n3283, S => n650, Z => n3285);
   U3818 : MUX2_X1 port map( A => REGISTERS_17_25_port, B => 
                           REGISTERS_19_25_port, S => n602, Z => n3286);
   U3819 : MUX2_X1 port map( A => REGISTERS_16_25_port, B => 
                           REGISTERS_18_25_port, S => n602, Z => n3287);
   U3820 : MUX2_X1 port map( A => n3287, B => n3286, S => n650, Z => n3288);
   U3821 : MUX2_X1 port map( A => n3288, B => n3285, S => n583, Z => n3289);
   U3822 : MUX2_X1 port map( A => n3289, B => n3282, S => r3013_A_3_port, Z => 
                           n3290);
   U3823 : MUX2_X1 port map( A => REGISTERS_13_25_port, B => 
                           REGISTERS_15_25_port, S => n602, Z => n3291);
   U3824 : MUX2_X1 port map( A => REGISTERS_12_25_port, B => 
                           REGISTERS_14_25_port, S => n602, Z => n3292);
   U3825 : MUX2_X1 port map( A => n3292, B => n3291, S => n650, Z => n3293);
   U3826 : MUX2_X1 port map( A => REGISTERS_9_25_port, B => 
                           REGISTERS_11_25_port, S => n602, Z => n3294);
   U3827 : MUX2_X1 port map( A => REGISTERS_8_25_port, B => 
                           REGISTERS_10_25_port, S => n602, Z => n3295);
   U3828 : MUX2_X1 port map( A => n3295, B => n3294, S => n650, Z => n3296);
   U3829 : MUX2_X1 port map( A => n3296, B => n3293, S => n583, Z => n3297);
   U3830 : MUX2_X1 port map( A => REGISTERS_5_25_port, B => REGISTERS_7_25_port
                           , S => n602, Z => n3298);
   U3831 : MUX2_X1 port map( A => REGISTERS_4_25_port, B => REGISTERS_6_25_port
                           , S => n602, Z => n3299);
   U3832 : MUX2_X1 port map( A => n3299, B => n3298, S => n650, Z => n3300);
   U3833 : MUX2_X1 port map( A => REGISTERS_1_25_port, B => REGISTERS_3_25_port
                           , S => n602, Z => n3301);
   U3834 : MUX2_X1 port map( A => REGISTERS_0_25_port, B => REGISTERS_2_25_port
                           , S => n602, Z => n3302);
   U3835 : MUX2_X1 port map( A => n3302, B => n3301, S => n650, Z => n3303);
   U3836 : MUX2_X1 port map( A => n3303, B => n3300, S => n583, Z => n3304);
   U3837 : MUX2_X1 port map( A => n3304, B => n3297, S => r3013_A_3_port, Z => 
                           n3305);
   U3838 : MUX2_X1 port map( A => n3305, B => n3290, S => r3013_A_4_port, Z => 
                           n3306);
   U3839 : MUX2_X1 port map( A => n3306, B => n3275, S => ADD_RD2_5_port, Z => 
                           N4501);
   U3840 : MUX2_X1 port map( A => REGISTERS_37_26_port, B => 
                           REGISTERS_39_26_port, S => n602, Z => n3307);
   U3841 : MUX2_X1 port map( A => REGISTERS_36_26_port, B => 
                           REGISTERS_38_26_port, S => n602, Z => n3308);
   U3842 : MUX2_X1 port map( A => n3308, B => n3307, S => n650, Z => n3309);
   U3843 : MUX2_X1 port map( A => REGISTERS_33_26_port, B => 
                           REGISTERS_35_26_port, S => n601, Z => n3310);
   U3844 : MUX2_X1 port map( A => REGISTERS_32_26_port, B => 
                           REGISTERS_34_26_port, S => n601, Z => n3311);
   U3845 : MUX2_X1 port map( A => n3311, B => n3310, S => n650, Z => n3312);
   U3846 : MUX2_X1 port map( A => n3312, B => n3309, S => n583, Z => n3313);
   U3847 : MUX2_X1 port map( A => REGISTERS_29_26_port, B => 
                           REGISTERS_31_26_port, S => n601, Z => n3314);
   U3848 : MUX2_X1 port map( A => REGISTERS_28_26_port, B => 
                           REGISTERS_30_26_port, S => n601, Z => n3315);
   U3849 : MUX2_X1 port map( A => n3315, B => n3314, S => n649, Z => n3316);
   U3850 : MUX2_X1 port map( A => REGISTERS_25_26_port, B => 
                           REGISTERS_27_26_port, S => n601, Z => n3317);
   U3851 : MUX2_X1 port map( A => REGISTERS_24_26_port, B => 
                           REGISTERS_26_26_port, S => n601, Z => n3318);
   U3852 : MUX2_X1 port map( A => n3318, B => n3317, S => n649, Z => n3319);
   U3853 : MUX2_X1 port map( A => n3319, B => n3316, S => n583, Z => n3320);
   U3854 : MUX2_X1 port map( A => REGISTERS_21_26_port, B => 
                           REGISTERS_23_26_port, S => n601, Z => n3321);
   U3855 : MUX2_X1 port map( A => REGISTERS_20_26_port, B => 
                           REGISTERS_22_26_port, S => n601, Z => n3322);
   U3856 : MUX2_X1 port map( A => n3322, B => n3321, S => n649, Z => n3323);
   U3857 : MUX2_X1 port map( A => REGISTERS_17_26_port, B => 
                           REGISTERS_19_26_port, S => n601, Z => n3324);
   U3858 : MUX2_X1 port map( A => REGISTERS_16_26_port, B => 
                           REGISTERS_18_26_port, S => n601, Z => n3325);
   U3859 : MUX2_X1 port map( A => n3325, B => n3324, S => n649, Z => n3326);
   U3860 : MUX2_X1 port map( A => n3326, B => n3323, S => n583, Z => n3327);
   U3861 : MUX2_X1 port map( A => n3327, B => n3320, S => r3013_A_3_port, Z => 
                           n3328);
   U3862 : MUX2_X1 port map( A => REGISTERS_13_26_port, B => 
                           REGISTERS_15_26_port, S => n601, Z => n3329);
   U3863 : MUX2_X1 port map( A => REGISTERS_12_26_port, B => 
                           REGISTERS_14_26_port, S => n601, Z => n3330);
   U3864 : MUX2_X1 port map( A => n3330, B => n3329, S => n649, Z => n3331);
   U3865 : MUX2_X1 port map( A => REGISTERS_9_26_port, B => 
                           REGISTERS_11_26_port, S => n601, Z => n3332);
   U3866 : MUX2_X1 port map( A => REGISTERS_8_26_port, B => 
                           REGISTERS_10_26_port, S => n601, Z => n3333);
   U3867 : MUX2_X1 port map( A => n3333, B => n3332, S => n649, Z => n3334);
   U3868 : MUX2_X1 port map( A => n3334, B => n3331, S => n583, Z => n3335);
   U3869 : MUX2_X1 port map( A => REGISTERS_5_26_port, B => REGISTERS_7_26_port
                           , S => n601, Z => n3336);
   U3870 : MUX2_X1 port map( A => REGISTERS_4_26_port, B => REGISTERS_6_26_port
                           , S => n600, Z => n3337);
   U3871 : MUX2_X1 port map( A => n3337, B => n3336, S => n649, Z => n3338);
   U3872 : MUX2_X1 port map( A => REGISTERS_1_26_port, B => REGISTERS_3_26_port
                           , S => n600, Z => n3339);
   U3873 : MUX2_X1 port map( A => REGISTERS_0_26_port, B => REGISTERS_2_26_port
                           , S => n600, Z => n3340);
   U3874 : MUX2_X1 port map( A => n3340, B => n3339, S => n649, Z => n3341);
   U3875 : MUX2_X1 port map( A => n3341, B => n3338, S => n583, Z => n3342);
   U3876 : MUX2_X1 port map( A => n3342, B => n3335, S => r3013_A_3_port, Z => 
                           n3343);
   U3877 : MUX2_X1 port map( A => n3343, B => n3328, S => r3013_A_4_port, Z => 
                           n3344);
   U3878 : MUX2_X1 port map( A => n3344, B => n3313, S => ADD_RD2_5_port, Z => 
                           N4500);
   U3879 : MUX2_X1 port map( A => REGISTERS_37_27_port, B => 
                           REGISTERS_39_27_port, S => n600, Z => n3345);
   U3880 : MUX2_X1 port map( A => REGISTERS_36_27_port, B => 
                           REGISTERS_38_27_port, S => n600, Z => n3346);
   U3881 : MUX2_X1 port map( A => n3346, B => n3345, S => n649, Z => n3347);
   U3882 : MUX2_X1 port map( A => REGISTERS_33_27_port, B => 
                           REGISTERS_35_27_port, S => n600, Z => n3348);
   U3883 : MUX2_X1 port map( A => REGISTERS_32_27_port, B => 
                           REGISTERS_34_27_port, S => n600, Z => n3349);
   U3884 : MUX2_X1 port map( A => n3349, B => n3348, S => n649, Z => n3350);
   U3885 : MUX2_X1 port map( A => n3350, B => n3347, S => n582, Z => n3351);
   U3886 : MUX2_X1 port map( A => REGISTERS_29_27_port, B => 
                           REGISTERS_31_27_port, S => n600, Z => n3352);
   U3887 : MUX2_X1 port map( A => REGISTERS_28_27_port, B => 
                           REGISTERS_30_27_port, S => n600, Z => n3353);
   U3888 : MUX2_X1 port map( A => n3353, B => n3352, S => n649, Z => n3354);
   U3889 : MUX2_X1 port map( A => REGISTERS_25_27_port, B => 
                           REGISTERS_27_27_port, S => n600, Z => n3355);
   U3890 : MUX2_X1 port map( A => REGISTERS_24_27_port, B => 
                           REGISTERS_26_27_port, S => n600, Z => n3356);
   U3891 : MUX2_X1 port map( A => n3356, B => n3355, S => n649, Z => n3357);
   U3892 : MUX2_X1 port map( A => n3357, B => n3354, S => n582, Z => n3358);
   U3893 : MUX2_X1 port map( A => REGISTERS_21_27_port, B => 
                           REGISTERS_23_27_port, S => n600, Z => n3359);
   U3894 : MUX2_X1 port map( A => REGISTERS_20_27_port, B => 
                           REGISTERS_22_27_port, S => n600, Z => n3360);
   U3895 : MUX2_X1 port map( A => n3360, B => n3359, S => n649, Z => n3361);
   U3896 : MUX2_X1 port map( A => REGISTERS_17_27_port, B => 
                           REGISTERS_19_27_port, S => n600, Z => n3362);
   U3897 : MUX2_X1 port map( A => REGISTERS_16_27_port, B => 
                           REGISTERS_18_27_port, S => n600, Z => n3363);
   U3898 : MUX2_X1 port map( A => n3363, B => n3362, S => n649, Z => n3364);
   U3899 : MUX2_X1 port map( A => n3364, B => n3361, S => n582, Z => n3365);
   U3900 : MUX2_X1 port map( A => n3365, B => n3358, S => r3013_A_3_port, Z => 
                           n3366);
   U3901 : MUX2_X1 port map( A => REGISTERS_13_27_port, B => 
                           REGISTERS_15_27_port, S => n599, Z => n3367);
   U3902 : MUX2_X1 port map( A => REGISTERS_12_27_port, B => 
                           REGISTERS_14_27_port, S => n599, Z => n3368);
   U3903 : MUX2_X1 port map( A => n3368, B => n3367, S => n649, Z => n3369);
   U3904 : MUX2_X1 port map( A => REGISTERS_9_27_port, B => 
                           REGISTERS_11_27_port, S => n599, Z => n3370);
   U3905 : MUX2_X1 port map( A => REGISTERS_8_27_port, B => 
                           REGISTERS_10_27_port, S => n599, Z => n3371);
   U3906 : MUX2_X1 port map( A => n3371, B => n3370, S => n648, Z => n3372);
   U3907 : MUX2_X1 port map( A => n3372, B => n3369, S => n582, Z => n3373);
   U3908 : MUX2_X1 port map( A => REGISTERS_5_27_port, B => REGISTERS_7_27_port
                           , S => n599, Z => n3374);
   U3909 : MUX2_X1 port map( A => REGISTERS_4_27_port, B => REGISTERS_6_27_port
                           , S => n599, Z => n3375);
   U3910 : MUX2_X1 port map( A => n3375, B => n3374, S => n648, Z => n3376);
   U3911 : MUX2_X1 port map( A => REGISTERS_1_27_port, B => REGISTERS_3_27_port
                           , S => n599, Z => n3377);
   U3912 : MUX2_X1 port map( A => REGISTERS_0_27_port, B => REGISTERS_2_27_port
                           , S => n599, Z => n3378);
   U3913 : MUX2_X1 port map( A => n3378, B => n3377, S => n648, Z => n3379);
   U3914 : MUX2_X1 port map( A => n3379, B => n3376, S => n582, Z => n3380);
   U3915 : MUX2_X1 port map( A => n3380, B => n3373, S => r3013_A_3_port, Z => 
                           n3381);
   U3916 : MUX2_X1 port map( A => n3381, B => n3366, S => r3013_A_4_port, Z => 
                           n3382);
   U3917 : MUX2_X1 port map( A => n3382, B => n3351, S => ADD_RD2_5_port, Z => 
                           N4499);
   U3918 : MUX2_X1 port map( A => REGISTERS_37_28_port, B => 
                           REGISTERS_39_28_port, S => n599, Z => n3383);
   U3919 : MUX2_X1 port map( A => REGISTERS_36_28_port, B => 
                           REGISTERS_38_28_port, S => n599, Z => n3384);
   U3920 : MUX2_X1 port map( A => n3384, B => n3383, S => n648, Z => n3385);
   U3921 : MUX2_X1 port map( A => REGISTERS_33_28_port, B => 
                           REGISTERS_35_28_port, S => n599, Z => n3386);
   U3922 : MUX2_X1 port map( A => REGISTERS_32_28_port, B => 
                           REGISTERS_34_28_port, S => n599, Z => n3387);
   U3923 : MUX2_X1 port map( A => n3387, B => n3386, S => n648, Z => n3388);
   U3924 : MUX2_X1 port map( A => n3388, B => n3385, S => n582, Z => n3389);
   U3925 : MUX2_X1 port map( A => REGISTERS_29_28_port, B => 
                           REGISTERS_31_28_port, S => n599, Z => n3390);
   U3926 : MUX2_X1 port map( A => REGISTERS_28_28_port, B => 
                           REGISTERS_30_28_port, S => n599, Z => n3391);
   U3927 : MUX2_X1 port map( A => n3391, B => n3390, S => n648, Z => n3392);
   U3928 : MUX2_X1 port map( A => REGISTERS_25_28_port, B => 
                           REGISTERS_27_28_port, S => n599, Z => n3393);
   U3929 : MUX2_X1 port map( A => REGISTERS_24_28_port, B => 
                           REGISTERS_26_28_port, S => n598, Z => n3394);
   U3930 : MUX2_X1 port map( A => n3394, B => n3393, S => n648, Z => n3395);
   U3931 : MUX2_X1 port map( A => n3395, B => n3392, S => n582, Z => n3396);
   U3932 : MUX2_X1 port map( A => REGISTERS_21_28_port, B => 
                           REGISTERS_23_28_port, S => n598, Z => n3397);
   U3933 : MUX2_X1 port map( A => REGISTERS_20_28_port, B => 
                           REGISTERS_22_28_port, S => n598, Z => n3398);
   U3934 : MUX2_X1 port map( A => n3398, B => n3397, S => n648, Z => n3399);
   U3935 : MUX2_X1 port map( A => REGISTERS_17_28_port, B => 
                           REGISTERS_19_28_port, S => n598, Z => n3400);
   U3936 : MUX2_X1 port map( A => REGISTERS_16_28_port, B => 
                           REGISTERS_18_28_port, S => n598, Z => n3401);
   U3937 : MUX2_X1 port map( A => n3401, B => n3400, S => n648, Z => n3402);
   U3938 : MUX2_X1 port map( A => n3402, B => n3399, S => n582, Z => n3403);
   U3939 : MUX2_X1 port map( A => n3403, B => n3396, S => r3013_A_3_port, Z => 
                           n3404);
   U3940 : MUX2_X1 port map( A => REGISTERS_13_28_port, B => 
                           REGISTERS_15_28_port, S => n598, Z => n3405);
   U3941 : MUX2_X1 port map( A => REGISTERS_12_28_port, B => 
                           REGISTERS_14_28_port, S => n598, Z => n3406);
   U3942 : MUX2_X1 port map( A => n3406, B => n3405, S => n648, Z => n3407);
   U3943 : MUX2_X1 port map( A => REGISTERS_9_28_port, B => 
                           REGISTERS_11_28_port, S => n598, Z => n3408);
   U3944 : MUX2_X1 port map( A => REGISTERS_8_28_port, B => 
                           REGISTERS_10_28_port, S => n598, Z => n3409);
   U3945 : MUX2_X1 port map( A => n3409, B => n3408, S => n648, Z => n3410);
   U3946 : MUX2_X1 port map( A => n3410, B => n3407, S => n582, Z => n3411);
   U3947 : MUX2_X1 port map( A => REGISTERS_5_28_port, B => REGISTERS_7_28_port
                           , S => n598, Z => n3412);
   U3948 : MUX2_X1 port map( A => REGISTERS_4_28_port, B => REGISTERS_6_28_port
                           , S => n598, Z => n3413);
   U3949 : MUX2_X1 port map( A => n3413, B => n3412, S => n648, Z => n3414);
   U3950 : MUX2_X1 port map( A => REGISTERS_1_28_port, B => REGISTERS_3_28_port
                           , S => n598, Z => n3415);
   U3951 : MUX2_X1 port map( A => REGISTERS_0_28_port, B => REGISTERS_2_28_port
                           , S => n598, Z => n3416);
   U3952 : MUX2_X1 port map( A => n3416, B => n3415, S => n648, Z => n3417);
   U3953 : MUX2_X1 port map( A => n3417, B => n3414, S => n582, Z => n3418);
   U3954 : MUX2_X1 port map( A => n3418, B => n3411, S => r3013_A_3_port, Z => 
                           n3419);
   U3955 : MUX2_X1 port map( A => n3419, B => n3404, S => r3013_A_4_port, Z => 
                           n3420);
   U3956 : MUX2_X1 port map( A => n3420, B => n3389, S => ADD_RD2_5_port, Z => 
                           N4498);
   U3957 : MUX2_X1 port map( A => REGISTERS_37_29_port, B => 
                           REGISTERS_39_29_port, S => n598, Z => n3421);
   U3958 : MUX2_X1 port map( A => REGISTERS_36_29_port, B => 
                           REGISTERS_38_29_port, S => n598, Z => n3422);
   U3959 : MUX2_X1 port map( A => n3422, B => n3421, S => n648, Z => n3423);
   U3960 : MUX2_X1 port map( A => REGISTERS_33_29_port, B => 
                           REGISTERS_35_29_port, S => n597, Z => n3424);
   U3961 : MUX2_X1 port map( A => REGISTERS_32_29_port, B => 
                           REGISTERS_34_29_port, S => n597, Z => n3425);
   U3962 : MUX2_X1 port map( A => n3425, B => n3424, S => n648, Z => n3426);
   U3963 : MUX2_X1 port map( A => n3426, B => n3423, S => n582, Z => n3427);
   U3964 : MUX2_X1 port map( A => REGISTERS_29_29_port, B => 
                           REGISTERS_31_29_port, S => n597, Z => n3428);
   U3965 : MUX2_X1 port map( A => REGISTERS_28_29_port, B => 
                           REGISTERS_30_29_port, S => n597, Z => n3429);
   U3966 : MUX2_X1 port map( A => n3429, B => n3428, S => n647, Z => n3430);
   U3967 : MUX2_X1 port map( A => REGISTERS_25_29_port, B => 
                           REGISTERS_27_29_port, S => n597, Z => n3431);
   U3968 : MUX2_X1 port map( A => REGISTERS_24_29_port, B => 
                           REGISTERS_26_29_port, S => n597, Z => n3432);
   U3969 : MUX2_X1 port map( A => n3432, B => n3431, S => n647, Z => n3433);
   U3970 : MUX2_X1 port map( A => n3433, B => n3430, S => n582, Z => n3434);
   U3971 : MUX2_X1 port map( A => REGISTERS_21_29_port, B => 
                           REGISTERS_23_29_port, S => n597, Z => n3435);
   U3972 : MUX2_X1 port map( A => REGISTERS_20_29_port, B => 
                           REGISTERS_22_29_port, S => n597, Z => n3436);
   U3973 : MUX2_X1 port map( A => n3436, B => n3435, S => n647, Z => n3437);
   U3974 : MUX2_X1 port map( A => REGISTERS_17_29_port, B => 
                           REGISTERS_19_29_port, S => n597, Z => n3438);
   U3975 : MUX2_X1 port map( A => REGISTERS_16_29_port, B => 
                           REGISTERS_18_29_port, S => n597, Z => n3439);
   U3976 : MUX2_X1 port map( A => n3439, B => n3438, S => n647, Z => n3440);
   U3977 : MUX2_X1 port map( A => n3440, B => n3437, S => n582, Z => n3441);
   U3978 : MUX2_X1 port map( A => n3441, B => n3434, S => r3013_A_3_port, Z => 
                           n3442);
   U3979 : MUX2_X1 port map( A => REGISTERS_13_29_port, B => 
                           REGISTERS_15_29_port, S => n597, Z => n3443);
   U3980 : MUX2_X1 port map( A => REGISTERS_12_29_port, B => 
                           REGISTERS_14_29_port, S => n597, Z => n3444);
   U3981 : MUX2_X1 port map( A => n3444, B => n3443, S => n647, Z => n3445);
   U3982 : MUX2_X1 port map( A => REGISTERS_9_29_port, B => 
                           REGISTERS_11_29_port, S => n597, Z => n3446);
   U3983 : MUX2_X1 port map( A => REGISTERS_8_29_port, B => 
                           REGISTERS_10_29_port, S => n597, Z => n3447);
   U3984 : MUX2_X1 port map( A => n3447, B => n3446, S => n647, Z => n3448);
   U3985 : MUX2_X1 port map( A => n3448, B => n3445, S => n581, Z => n3449);
   U3986 : MUX2_X1 port map( A => REGISTERS_5_29_port, B => REGISTERS_7_29_port
                           , S => n597, Z => n3450);
   U3987 : MUX2_X1 port map( A => REGISTERS_4_29_port, B => REGISTERS_6_29_port
                           , S => n596, Z => n3451);
   U3988 : MUX2_X1 port map( A => n3451, B => n3450, S => n647, Z => n3452);
   U3989 : MUX2_X1 port map( A => REGISTERS_1_29_port, B => REGISTERS_3_29_port
                           , S => n596, Z => n3453);
   U3990 : MUX2_X1 port map( A => REGISTERS_0_29_port, B => REGISTERS_2_29_port
                           , S => n596, Z => n3454);
   U3991 : MUX2_X1 port map( A => n3454, B => n3453, S => n647, Z => n3455);
   U3992 : MUX2_X1 port map( A => n3455, B => n3452, S => n581, Z => n3456);
   U3993 : MUX2_X1 port map( A => n3456, B => n3449, S => r3013_A_3_port, Z => 
                           n3457);
   U3994 : MUX2_X1 port map( A => n3457, B => n3442, S => r3013_A_4_port, Z => 
                           n3458);
   U3995 : MUX2_X1 port map( A => n3458, B => n3427, S => ADD_RD2_5_port, Z => 
                           N4497);
   U3996 : MUX2_X1 port map( A => REGISTERS_37_30_port, B => 
                           REGISTERS_39_30_port, S => n596, Z => n3459);
   U3997 : MUX2_X1 port map( A => REGISTERS_36_30_port, B => 
                           REGISTERS_38_30_port, S => n596, Z => n3460);
   U3998 : MUX2_X1 port map( A => n3460, B => n3459, S => n647, Z => n3461);
   U3999 : MUX2_X1 port map( A => REGISTERS_33_30_port, B => 
                           REGISTERS_35_30_port, S => n596, Z => n3462);
   U4000 : MUX2_X1 port map( A => REGISTERS_32_30_port, B => 
                           REGISTERS_34_30_port, S => n596, Z => n3463);
   U4001 : MUX2_X1 port map( A => n3463, B => n3462, S => n647, Z => n3464);
   U4002 : MUX2_X1 port map( A => n3464, B => n3461, S => n581, Z => n3465);
   U4003 : MUX2_X1 port map( A => REGISTERS_29_30_port, B => 
                           REGISTERS_31_30_port, S => n596, Z => n3466);
   U4004 : MUX2_X1 port map( A => REGISTERS_28_30_port, B => 
                           REGISTERS_30_30_port, S => n596, Z => n3467);
   U4005 : MUX2_X1 port map( A => n3467, B => n3466, S => n647, Z => n3468);
   U4006 : MUX2_X1 port map( A => REGISTERS_25_30_port, B => 
                           REGISTERS_27_30_port, S => n596, Z => n3469);
   U4007 : MUX2_X1 port map( A => REGISTERS_24_30_port, B => 
                           REGISTERS_26_30_port, S => n596, Z => n3470);
   U4008 : MUX2_X1 port map( A => n3470, B => n3469, S => n647, Z => n3471);
   U4009 : MUX2_X1 port map( A => n3471, B => n3468, S => n581, Z => n3472);
   U4010 : MUX2_X1 port map( A => REGISTERS_21_30_port, B => 
                           REGISTERS_23_30_port, S => n596, Z => n3473);
   U4011 : MUX2_X1 port map( A => REGISTERS_20_30_port, B => 
                           REGISTERS_22_30_port, S => n596, Z => n3474);
   U4012 : MUX2_X1 port map( A => n3474, B => n3473, S => n647, Z => n3475);
   U4013 : MUX2_X1 port map( A => REGISTERS_17_30_port, B => 
                           REGISTERS_19_30_port, S => n596, Z => n3476);
   U4014 : MUX2_X1 port map( A => REGISTERS_16_30_port, B => 
                           REGISTERS_18_30_port, S => n596, Z => n3477);
   U4015 : MUX2_X1 port map( A => n3477, B => n3476, S => n647, Z => n3478);
   U4016 : MUX2_X1 port map( A => n3478, B => n3475, S => n581, Z => n3479);
   U4017 : MUX2_X1 port map( A => n3479, B => n3472, S => r3013_A_3_port, Z => 
                           n3480);
   U4018 : MUX2_X1 port map( A => REGISTERS_13_30_port, B => 
                           REGISTERS_15_30_port, S => n595, Z => n3481);
   U4019 : MUX2_X1 port map( A => REGISTERS_12_30_port, B => 
                           REGISTERS_14_30_port, S => n595, Z => n3482);
   U4020 : MUX2_X1 port map( A => n3482, B => n3481, S => n647, Z => n3483);
   U4021 : MUX2_X1 port map( A => REGISTERS_9_30_port, B => 
                           REGISTERS_11_30_port, S => n595, Z => n3484);
   U4022 : MUX2_X1 port map( A => REGISTERS_8_30_port, B => 
                           REGISTERS_10_30_port, S => n595, Z => n3485);
   U4023 : MUX2_X1 port map( A => n3485, B => n3484, S => n646, Z => n3486);
   U4024 : MUX2_X1 port map( A => n3486, B => n3483, S => n581, Z => n3487);
   U4025 : MUX2_X1 port map( A => REGISTERS_5_30_port, B => REGISTERS_7_30_port
                           , S => n595, Z => n3488);
   U4026 : MUX2_X1 port map( A => REGISTERS_4_30_port, B => REGISTERS_6_30_port
                           , S => n595, Z => n3489);
   U4027 : MUX2_X1 port map( A => n3489, B => n3488, S => n646, Z => n3490);
   U4028 : MUX2_X1 port map( A => REGISTERS_1_30_port, B => REGISTERS_3_30_port
                           , S => n595, Z => n3491);
   U4029 : MUX2_X1 port map( A => REGISTERS_0_30_port, B => REGISTERS_2_30_port
                           , S => n595, Z => n3492);
   U4030 : MUX2_X1 port map( A => n3492, B => n3491, S => n646, Z => n3493);
   U4031 : MUX2_X1 port map( A => n3493, B => n3490, S => n581, Z => n3494);
   U4032 : MUX2_X1 port map( A => n3494, B => n3487, S => r3013_A_3_port, Z => 
                           n3495);
   U4033 : MUX2_X1 port map( A => n3495, B => n3480, S => r3013_A_4_port, Z => 
                           n3496);
   U4034 : MUX2_X1 port map( A => n3496, B => n3465, S => ADD_RD2_5_port, Z => 
                           N4496);
   U4035 : MUX2_X1 port map( A => REGISTERS_37_31_port, B => 
                           REGISTERS_39_31_port, S => n595, Z => n3497);
   U4036 : MUX2_X1 port map( A => REGISTERS_36_31_port, B => 
                           REGISTERS_38_31_port, S => n595, Z => n3498);
   U4037 : MUX2_X1 port map( A => n3498, B => n3497, S => n646, Z => n3499);
   U4038 : MUX2_X1 port map( A => REGISTERS_33_31_port, B => 
                           REGISTERS_35_31_port, S => n595, Z => n3500);
   U4039 : MUX2_X1 port map( A => REGISTERS_32_31_port, B => 
                           REGISTERS_34_31_port, S => n595, Z => n3501);
   U4040 : MUX2_X1 port map( A => n3501, B => n3500, S => n646, Z => n3502);
   U4041 : MUX2_X1 port map( A => n3502, B => n3499, S => n581, Z => n3503);
   U4042 : MUX2_X1 port map( A => REGISTERS_29_31_port, B => 
                           REGISTERS_31_31_port, S => n595, Z => n3504);
   U4043 : MUX2_X1 port map( A => REGISTERS_28_31_port, B => 
                           REGISTERS_30_31_port, S => n595, Z => n3505);
   U4044 : MUX2_X1 port map( A => n3505, B => n3504, S => n646, Z => n3506);
   U4045 : MUX2_X1 port map( A => REGISTERS_25_31_port, B => 
                           REGISTERS_27_31_port, S => n595, Z => n3507);
   U4046 : MUX2_X1 port map( A => REGISTERS_24_31_port, B => 
                           REGISTERS_26_31_port, S => n594, Z => n3508);
   U4047 : MUX2_X1 port map( A => n3508, B => n3507, S => n646, Z => n3509);
   U4048 : MUX2_X1 port map( A => n3509, B => n3506, S => n581, Z => n3510);
   U4049 : MUX2_X1 port map( A => REGISTERS_21_31_port, B => 
                           REGISTERS_23_31_port, S => n594, Z => n3511);
   U4050 : MUX2_X1 port map( A => REGISTERS_20_31_port, B => 
                           REGISTERS_22_31_port, S => n594, Z => n3512);
   U4051 : MUX2_X1 port map( A => n3512, B => n3511, S => n646, Z => n3513);
   U4052 : MUX2_X1 port map( A => REGISTERS_17_31_port, B => 
                           REGISTERS_19_31_port, S => n594, Z => n3514);
   U4053 : MUX2_X1 port map( A => REGISTERS_16_31_port, B => 
                           REGISTERS_18_31_port, S => n594, Z => n3515);
   U4054 : MUX2_X1 port map( A => n3515, B => n3514, S => n646, Z => n3516);
   U4055 : MUX2_X1 port map( A => n3516, B => n3513, S => n581, Z => n3517);
   U4056 : MUX2_X1 port map( A => n3517, B => n3510, S => r3013_A_3_port, Z => 
                           n3518);
   U4057 : MUX2_X1 port map( A => REGISTERS_13_31_port, B => 
                           REGISTERS_15_31_port, S => n594, Z => n3519);
   U4058 : MUX2_X1 port map( A => REGISTERS_12_31_port, B => 
                           REGISTERS_14_31_port, S => n594, Z => n3520);
   U4059 : MUX2_X1 port map( A => n3520, B => n3519, S => n646, Z => n3521);
   U4060 : MUX2_X1 port map( A => REGISTERS_9_31_port, B => 
                           REGISTERS_11_31_port, S => n594, Z => n3522);
   U4061 : MUX2_X1 port map( A => REGISTERS_8_31_port, B => 
                           REGISTERS_10_31_port, S => n594, Z => n3523);
   U4062 : MUX2_X1 port map( A => n3523, B => n3522, S => n646, Z => n3524);
   U4063 : MUX2_X1 port map( A => n3524, B => n3521, S => n581, Z => n3525);
   U4064 : MUX2_X1 port map( A => REGISTERS_5_31_port, B => REGISTERS_7_31_port
                           , S => n594, Z => n3526);
   U4065 : MUX2_X1 port map( A => REGISTERS_4_31_port, B => REGISTERS_6_31_port
                           , S => n594, Z => n3527);
   U4066 : MUX2_X1 port map( A => n3527, B => n3526, S => n646, Z => n3528);
   U4067 : MUX2_X1 port map( A => REGISTERS_1_31_port, B => REGISTERS_3_31_port
                           , S => n594, Z => n3529);
   U4068 : MUX2_X1 port map( A => REGISTERS_0_31_port, B => REGISTERS_2_31_port
                           , S => n594, Z => n3530);
   U4069 : MUX2_X1 port map( A => n3530, B => n3529, S => n646, Z => n3531);
   U4070 : MUX2_X1 port map( A => n3531, B => n3528, S => n581, Z => n3532);
   U4071 : MUX2_X1 port map( A => n3532, B => n3525, S => r3013_A_3_port, Z => 
                           n3533);
   U4072 : MUX2_X1 port map( A => n3533, B => n3518, S => r3013_A_4_port, Z => 
                           n3534);
   U4073 : MUX2_X1 port map( A => n3534, B => n3503, S => ADD_RD2_5_port, Z => 
                           N4495);
   U4074 : MUX2_X1 port map( A => REGISTERS_37_0_port, B => REGISTERS_39_0_port
                           , S => n722, Z => n3535);
   U4075 : MUX2_X1 port map( A => REGISTERS_36_0_port, B => REGISTERS_38_0_port
                           , S => n722, Z => n3536);
   U4076 : MUX2_X1 port map( A => n3536, B => n3535, S => n753, Z => n3537);
   U4077 : MUX2_X1 port map( A => REGISTERS_33_0_port, B => REGISTERS_35_0_port
                           , S => n722, Z => n3538);
   U4078 : MUX2_X1 port map( A => REGISTERS_32_0_port, B => REGISTERS_34_0_port
                           , S => n722, Z => n3539);
   U4079 : MUX2_X1 port map( A => n3539, B => n3538, S => n753, Z => n3540);
   U4080 : MUX2_X1 port map( A => n3540, B => n3537, S => n679, Z => n3541);
   U4081 : MUX2_X1 port map( A => REGISTERS_29_0_port, B => REGISTERS_31_0_port
                           , S => n722, Z => n3542);
   U4082 : MUX2_X1 port map( A => REGISTERS_28_0_port, B => REGISTERS_30_0_port
                           , S => n722, Z => n3543);
   U4083 : MUX2_X1 port map( A => n3543, B => n3542, S => n753, Z => n3544);
   U4084 : MUX2_X1 port map( A => REGISTERS_25_0_port, B => REGISTERS_27_0_port
                           , S => n722, Z => n3545);
   U4085 : MUX2_X1 port map( A => REGISTERS_24_0_port, B => REGISTERS_26_0_port
                           , S => n722, Z => n3546);
   U4086 : MUX2_X1 port map( A => n3546, B => n3545, S => n753, Z => n3547);
   U4087 : MUX2_X1 port map( A => n3547, B => n3544, S => n679, Z => n3548);
   U4088 : MUX2_X1 port map( A => REGISTERS_21_0_port, B => REGISTERS_23_0_port
                           , S => n722, Z => n3549);
   U4089 : MUX2_X1 port map( A => REGISTERS_20_0_port, B => REGISTERS_22_0_port
                           , S => n722, Z => n3550);
   U4090 : MUX2_X1 port map( A => n3550, B => n3549, S => n753, Z => n3551);
   U4091 : MUX2_X1 port map( A => REGISTERS_17_0_port, B => REGISTERS_19_0_port
                           , S => n722, Z => n3552);
   U4092 : MUX2_X1 port map( A => REGISTERS_16_0_port, B => REGISTERS_18_0_port
                           , S => n722, Z => n3553);
   U4093 : MUX2_X1 port map( A => n3553, B => n3552, S => n753, Z => n3554);
   U4094 : MUX2_X1 port map( A => n3554, B => n3551, S => n679, Z => n3555);
   U4095 : MUX2_X1 port map( A => n3555, B => n3548, S => r3007_A_3_port, Z => 
                           n3556);
   U4096 : MUX2_X1 port map( A => REGISTERS_13_0_port, B => REGISTERS_15_0_port
                           , S => n721, Z => n3557);
   U4097 : MUX2_X1 port map( A => REGISTERS_12_0_port, B => REGISTERS_14_0_port
                           , S => n721, Z => n3558);
   U4098 : MUX2_X1 port map( A => n3558, B => n3557, S => n753, Z => n3559);
   U4099 : MUX2_X1 port map( A => REGISTERS_9_0_port, B => REGISTERS_11_0_port,
                           S => n721, Z => n3560);
   U4100 : MUX2_X1 port map( A => REGISTERS_8_0_port, B => REGISTERS_10_0_port,
                           S => n721, Z => n3561);
   U4101 : MUX2_X1 port map( A => n3561, B => n3560, S => n752, Z => n3562);
   U4102 : MUX2_X1 port map( A => n3562, B => n3559, S => n679, Z => n3563);
   U4103 : MUX2_X1 port map( A => REGISTERS_5_0_port, B => REGISTERS_7_0_port, 
                           S => n721, Z => n3564_port);
   U4104 : MUX2_X1 port map( A => REGISTERS_4_0_port, B => REGISTERS_6_0_port, 
                           S => n721, Z => n3565_port);
   U4105 : MUX2_X1 port map( A => n3565_port, B => n3564_port, S => n752, Z => 
                           n3566_port);
   U4106 : MUX2_X1 port map( A => REGISTERS_1_0_port, B => REGISTERS_3_0_port, 
                           S => n721, Z => n3567_port);
   U4107 : MUX2_X1 port map( A => REGISTERS_0_0_port, B => REGISTERS_2_0_port, 
                           S => n721, Z => n3568_port);
   U4108 : MUX2_X1 port map( A => n3568_port, B => n3567_port, S => n752, Z => 
                           n3569_port);
   U4109 : MUX2_X1 port map( A => n3569_port, B => n3566_port, S => n679, Z => 
                           n3570_port);
   U4110 : MUX2_X1 port map( A => n3570_port, B => n3563, S => r3007_A_3_port, 
                           Z => n3571_port);
   U4111 : MUX2_X1 port map( A => n3571_port, B => n3556, S => r3007_A_4_port, 
                           Z => n3572_port);
   U4112 : MUX2_X1 port map( A => n3572_port, B => n3541, S => ADD_RD1_5_port, 
                           Z => N4420);
   U4113 : MUX2_X1 port map( A => REGISTERS_37_1_port, B => REGISTERS_39_1_port
                           , S => n721, Z => n3573);
   U4114 : MUX2_X1 port map( A => REGISTERS_36_1_port, B => REGISTERS_38_1_port
                           , S => n721, Z => n3574);
   U4115 : MUX2_X1 port map( A => n3574, B => n3573, S => n752, Z => n3575);
   U4116 : MUX2_X1 port map( A => REGISTERS_33_1_port, B => REGISTERS_35_1_port
                           , S => n721, Z => n3576);
   U4117 : MUX2_X1 port map( A => REGISTERS_32_1_port, B => REGISTERS_34_1_port
                           , S => n721, Z => n3577_port);
   U4118 : MUX2_X1 port map( A => n3577_port, B => n3576, S => n752, Z => 
                           n3578_port);
   U4119 : MUX2_X1 port map( A => n3578_port, B => n3575, S => n679, Z => 
                           n3579_port);
   U4120 : MUX2_X1 port map( A => REGISTERS_29_1_port, B => REGISTERS_31_1_port
                           , S => n721, Z => n3580_port);
   U4121 : MUX2_X1 port map( A => REGISTERS_28_1_port, B => REGISTERS_30_1_port
                           , S => n721, Z => n3581_port);
   U4122 : MUX2_X1 port map( A => n3581_port, B => n3580_port, S => n752, Z => 
                           n3582_port);
   U4123 : MUX2_X1 port map( A => REGISTERS_25_1_port, B => REGISTERS_27_1_port
                           , S => n721, Z => n3583_port);
   U4124 : MUX2_X1 port map( A => REGISTERS_24_1_port, B => REGISTERS_26_1_port
                           , S => n720, Z => n3584_port);
   U4125 : MUX2_X1 port map( A => n3584_port, B => n3583_port, S => n752, Z => 
                           n3585_port);
   U4126 : MUX2_X1 port map( A => n3585_port, B => n3582_port, S => n679, Z => 
                           n3586);
   U4127 : MUX2_X1 port map( A => REGISTERS_21_1_port, B => REGISTERS_23_1_port
                           , S => n720, Z => n3587);
   U4128 : MUX2_X1 port map( A => REGISTERS_20_1_port, B => REGISTERS_22_1_port
                           , S => n720, Z => n3588);
   U4129 : MUX2_X1 port map( A => n3588, B => n3587, S => n752, Z => n3589);
   U4130 : MUX2_X1 port map( A => REGISTERS_17_1_port, B => REGISTERS_19_1_port
                           , S => n720, Z => n3590_port);
   U4131 : MUX2_X1 port map( A => REGISTERS_16_1_port, B => REGISTERS_18_1_port
                           , S => n720, Z => n3591_port);
   U4132 : MUX2_X1 port map( A => n3591_port, B => n3590_port, S => n752, Z => 
                           n3592_port);
   U4133 : MUX2_X1 port map( A => n3592_port, B => n3589, S => n678, Z => 
                           n3593_port);
   U4134 : MUX2_X1 port map( A => n3593_port, B => n3586, S => r3007_A_3_port, 
                           Z => n3594_port);
   U4135 : MUX2_X1 port map( A => REGISTERS_13_1_port, B => REGISTERS_15_1_port
                           , S => n720, Z => n3595_port);
   U4136 : MUX2_X1 port map( A => REGISTERS_12_1_port, B => REGISTERS_14_1_port
                           , S => n720, Z => n3596_port);
   U4137 : MUX2_X1 port map( A => n3596_port, B => n3595_port, S => n752, Z => 
                           n3597_port);
   U4138 : MUX2_X1 port map( A => REGISTERS_9_1_port, B => REGISTERS_11_1_port,
                           S => n720, Z => n3598_port);
   U4139 : MUX2_X1 port map( A => REGISTERS_8_1_port, B => REGISTERS_10_1_port,
                           S => n720, Z => n3599);
   U4140 : MUX2_X1 port map( A => n3599, B => n3598_port, S => n752, Z => n3600
                           );
   U4141 : MUX2_X1 port map( A => n3600, B => n3597_port, S => n678, Z => n3601
                           );
   U4142 : MUX2_X1 port map( A => REGISTERS_5_1_port, B => REGISTERS_7_1_port, 
                           S => n720, Z => n3602);
   U4143 : MUX2_X1 port map( A => REGISTERS_4_1_port, B => REGISTERS_6_1_port, 
                           S => n720, Z => n3603);
   U4144 : MUX2_X1 port map( A => n3603, B => n3602, S => n752, Z => n3604);
   U4145 : MUX2_X1 port map( A => REGISTERS_1_1_port, B => REGISTERS_3_1_port, 
                           S => n720, Z => n3605);
   U4146 : MUX2_X1 port map( A => REGISTERS_0_1_port, B => REGISTERS_2_1_port, 
                           S => n720, Z => n3606);
   U4147 : MUX2_X1 port map( A => n3606, B => n3605, S => n752, Z => n3607);
   U4148 : MUX2_X1 port map( A => n3607, B => n3604, S => n678, Z => n3608);
   U4149 : MUX2_X1 port map( A => n3608, B => n3601, S => r3007_A_3_port, Z => 
                           n3609);
   U4150 : MUX2_X1 port map( A => n3609, B => n3594_port, S => r3007_A_4_port, 
                           Z => n3610);
   U4151 : MUX2_X1 port map( A => n3610, B => n3579_port, S => ADD_RD1_5_port, 
                           Z => N4419);
   U4152 : MUX2_X1 port map( A => REGISTERS_37_2_port, B => REGISTERS_39_2_port
                           , S => n720, Z => n3611);
   U4153 : MUX2_X1 port map( A => REGISTERS_36_2_port, B => REGISTERS_38_2_port
                           , S => n720, Z => n3612);
   U4154 : MUX2_X1 port map( A => n3612, B => n3611, S => n752, Z => n3613);
   U4155 : MUX2_X1 port map( A => REGISTERS_33_2_port, B => REGISTERS_35_2_port
                           , S => n719, Z => n3614);
   U4156 : MUX2_X1 port map( A => REGISTERS_32_2_port, B => REGISTERS_34_2_port
                           , S => n719, Z => n3615);
   U4157 : MUX2_X1 port map( A => n3615, B => n3614, S => n752, Z => n3616);
   U4158 : MUX2_X1 port map( A => n3616, B => n3613, S => n678, Z => n3617);
   U4159 : MUX2_X1 port map( A => REGISTERS_29_2_port, B => REGISTERS_31_2_port
                           , S => n719, Z => n3618);
   U4160 : MUX2_X1 port map( A => REGISTERS_28_2_port, B => REGISTERS_30_2_port
                           , S => n719, Z => n3619);
   U4161 : MUX2_X1 port map( A => n3619, B => n3618, S => n751, Z => n3620);
   U4162 : MUX2_X1 port map( A => REGISTERS_25_2_port, B => REGISTERS_27_2_port
                           , S => n719, Z => n3621);
   U4163 : MUX2_X1 port map( A => REGISTERS_24_2_port, B => REGISTERS_26_2_port
                           , S => n719, Z => n3622);
   U4164 : MUX2_X1 port map( A => n3622, B => n3621, S => n751, Z => n3623);
   U4165 : MUX2_X1 port map( A => n3623, B => n3620, S => n678, Z => n3624);
   U4166 : MUX2_X1 port map( A => REGISTERS_21_2_port, B => REGISTERS_23_2_port
                           , S => n719, Z => n3625);
   U4167 : MUX2_X1 port map( A => REGISTERS_20_2_port, B => REGISTERS_22_2_port
                           , S => n719, Z => n3626);
   U4168 : MUX2_X1 port map( A => n3626, B => n3625, S => n751, Z => n3627);
   U4169 : MUX2_X1 port map( A => REGISTERS_17_2_port, B => REGISTERS_19_2_port
                           , S => n719, Z => n3628);
   U4170 : MUX2_X1 port map( A => REGISTERS_16_2_port, B => REGISTERS_18_2_port
                           , S => n719, Z => n3629);
   U4171 : MUX2_X1 port map( A => n3629, B => n3628, S => n751, Z => n3630);
   U4172 : MUX2_X1 port map( A => n3630, B => n3627, S => n678, Z => n3631);
   U4173 : MUX2_X1 port map( A => n3631, B => n3624, S => r3007_A_3_port, Z => 
                           n3632);
   U4174 : MUX2_X1 port map( A => REGISTERS_13_2_port, B => REGISTERS_15_2_port
                           , S => n719, Z => n3633);
   U4175 : MUX2_X1 port map( A => REGISTERS_12_2_port, B => REGISTERS_14_2_port
                           , S => n719, Z => n3634);
   U4176 : MUX2_X1 port map( A => n3634, B => n3633, S => n751, Z => n3635);
   U4177 : MUX2_X1 port map( A => REGISTERS_9_2_port, B => REGISTERS_11_2_port,
                           S => n719, Z => n3636);
   U4178 : MUX2_X1 port map( A => REGISTERS_8_2_port, B => REGISTERS_10_2_port,
                           S => n719, Z => n3637);
   U4179 : MUX2_X1 port map( A => n3637, B => n3636, S => n751, Z => n3638);
   U4180 : MUX2_X1 port map( A => n3638, B => n3635, S => n678, Z => n3639);
   U4181 : MUX2_X1 port map( A => REGISTERS_5_2_port, B => REGISTERS_7_2_port, 
                           S => n719, Z => n3640);
   U4182 : MUX2_X1 port map( A => REGISTERS_4_2_port, B => REGISTERS_6_2_port, 
                           S => n718, Z => n3641);
   U4183 : MUX2_X1 port map( A => n3641, B => n3640, S => n751, Z => n3642);
   U4184 : MUX2_X1 port map( A => REGISTERS_1_2_port, B => REGISTERS_3_2_port, 
                           S => n718, Z => n3643);
   U4185 : MUX2_X1 port map( A => REGISTERS_0_2_port, B => REGISTERS_2_2_port, 
                           S => n718, Z => n3644);
   U4186 : MUX2_X1 port map( A => n3644, B => n3643, S => n751, Z => n3645);
   U4187 : MUX2_X1 port map( A => n3645, B => n3642, S => n678, Z => n3646);
   U4188 : MUX2_X1 port map( A => n3646, B => n3639, S => r3007_A_3_port, Z => 
                           n3647);
   U4189 : MUX2_X1 port map( A => n3647, B => n3632, S => r3007_A_4_port, Z => 
                           n3648);
   U4190 : MUX2_X1 port map( A => n3648, B => n3617, S => ADD_RD1_5_port, Z => 
                           N4418);
   U4191 : MUX2_X1 port map( A => REGISTERS_37_3_port, B => REGISTERS_39_3_port
                           , S => n718, Z => n3649);
   U4192 : MUX2_X1 port map( A => REGISTERS_36_3_port, B => REGISTERS_38_3_port
                           , S => n718, Z => n3650);
   U4193 : MUX2_X1 port map( A => n3650, B => n3649, S => n751, Z => n3651);
   U4194 : MUX2_X1 port map( A => REGISTERS_33_3_port, B => REGISTERS_35_3_port
                           , S => n718, Z => n3652);
   U4195 : MUX2_X1 port map( A => REGISTERS_32_3_port, B => REGISTERS_34_3_port
                           , S => n718, Z => n3653);
   U4196 : MUX2_X1 port map( A => n3653, B => n3652, S => n751, Z => n3654);
   U4197 : MUX2_X1 port map( A => n3654, B => n3651, S => n678, Z => n3655);
   U4198 : MUX2_X1 port map( A => REGISTERS_29_3_port, B => REGISTERS_31_3_port
                           , S => n718, Z => n3656);
   U4199 : MUX2_X1 port map( A => REGISTERS_28_3_port, B => REGISTERS_30_3_port
                           , S => n718, Z => n3657);
   U4200 : MUX2_X1 port map( A => n3657, B => n3656, S => n751, Z => n3658);
   U4201 : MUX2_X1 port map( A => REGISTERS_25_3_port, B => REGISTERS_27_3_port
                           , S => n718, Z => n3659);
   U4202 : MUX2_X1 port map( A => REGISTERS_24_3_port, B => REGISTERS_26_3_port
                           , S => n718, Z => n3660);
   U4203 : MUX2_X1 port map( A => n3660, B => n3659, S => n751, Z => n3661);
   U4204 : MUX2_X1 port map( A => n3661, B => n3658, S => n678, Z => n3662);
   U4205 : MUX2_X1 port map( A => REGISTERS_21_3_port, B => REGISTERS_23_3_port
                           , S => n718, Z => n3663);
   U4206 : MUX2_X1 port map( A => REGISTERS_20_3_port, B => REGISTERS_22_3_port
                           , S => n718, Z => n3664);
   U4207 : MUX2_X1 port map( A => n3664, B => n3663, S => n751, Z => n3665);
   U4208 : MUX2_X1 port map( A => REGISTERS_17_3_port, B => REGISTERS_19_3_port
                           , S => n718, Z => n3666);
   U4209 : MUX2_X1 port map( A => REGISTERS_16_3_port, B => REGISTERS_18_3_port
                           , S => n718, Z => n3667);
   U4210 : MUX2_X1 port map( A => n3667, B => n3666, S => n751, Z => n3668);
   U4211 : MUX2_X1 port map( A => n3668, B => n3665, S => n678, Z => n3669);
   U4212 : MUX2_X1 port map( A => n3669, B => n3662, S => r3007_A_3_port, Z => 
                           n3670);
   U4213 : MUX2_X1 port map( A => REGISTERS_13_3_port, B => REGISTERS_15_3_port
                           , S => n717, Z => n3671);
   U4214 : MUX2_X1 port map( A => REGISTERS_12_3_port, B => REGISTERS_14_3_port
                           , S => n717, Z => n3672);
   U4215 : MUX2_X1 port map( A => n3672, B => n3671, S => n751, Z => n3673);
   U4216 : MUX2_X1 port map( A => REGISTERS_9_3_port, B => REGISTERS_11_3_port,
                           S => n717, Z => n3674);
   U4217 : MUX2_X1 port map( A => REGISTERS_8_3_port, B => REGISTERS_10_3_port,
                           S => n717, Z => n3675);
   U4218 : MUX2_X1 port map( A => n3675, B => n3674, S => n750, Z => n3676);
   U4219 : MUX2_X1 port map( A => n3676, B => n3673, S => n678, Z => n3677);
   U4220 : MUX2_X1 port map( A => REGISTERS_5_3_port, B => REGISTERS_7_3_port, 
                           S => n717, Z => n3678);
   U4221 : MUX2_X1 port map( A => REGISTERS_4_3_port, B => REGISTERS_6_3_port, 
                           S => n717, Z => n3679);
   U4222 : MUX2_X1 port map( A => n3679, B => n3678, S => n750, Z => n3680);
   U4223 : MUX2_X1 port map( A => REGISTERS_1_3_port, B => REGISTERS_3_3_port, 
                           S => n717, Z => n3681);
   U4224 : MUX2_X1 port map( A => REGISTERS_0_3_port, B => REGISTERS_2_3_port, 
                           S => n717, Z => n3682);
   U4225 : MUX2_X1 port map( A => n3682, B => n3681, S => n750, Z => n3683);
   U4226 : MUX2_X1 port map( A => n3683, B => n3680, S => n678, Z => n3684);
   U4227 : MUX2_X1 port map( A => n3684, B => n3677, S => r3007_A_3_port, Z => 
                           n3685);
   U4228 : MUX2_X1 port map( A => n3685, B => n3670, S => r3007_A_4_port, Z => 
                           n3686);
   U4229 : MUX2_X1 port map( A => n3686, B => n3655, S => ADD_RD1_5_port, Z => 
                           N4417);
   U4230 : MUX2_X1 port map( A => REGISTERS_37_4_port, B => REGISTERS_39_4_port
                           , S => n717, Z => n3687);
   U4231 : MUX2_X1 port map( A => REGISTERS_36_4_port, B => REGISTERS_38_4_port
                           , S => n717, Z => n3688);
   U4232 : MUX2_X1 port map( A => n3688, B => n3687, S => n750, Z => n3689);
   U4233 : MUX2_X1 port map( A => REGISTERS_33_4_port, B => REGISTERS_35_4_port
                           , S => n717, Z => n3690);
   U4234 : MUX2_X1 port map( A => REGISTERS_32_4_port, B => REGISTERS_34_4_port
                           , S => n717, Z => n3691);
   U4235 : MUX2_X1 port map( A => n3691, B => n3690, S => n750, Z => n3692);
   U4236 : MUX2_X1 port map( A => n3692, B => n3689, S => n678, Z => n3693);
   U4237 : MUX2_X1 port map( A => REGISTERS_29_4_port, B => REGISTERS_31_4_port
                           , S => n717, Z => n3694);
   U4238 : MUX2_X1 port map( A => REGISTERS_28_4_port, B => REGISTERS_30_4_port
                           , S => n717, Z => n3695);
   U4239 : MUX2_X1 port map( A => n3695, B => n3694, S => n750, Z => n3696);
   U4240 : MUX2_X1 port map( A => REGISTERS_25_4_port, B => REGISTERS_27_4_port
                           , S => n717, Z => n3697);
   U4241 : MUX2_X1 port map( A => REGISTERS_24_4_port, B => REGISTERS_26_4_port
                           , S => n716, Z => n3698);
   U4242 : MUX2_X1 port map( A => n3698, B => n3697, S => n750, Z => n3699);
   U4243 : MUX2_X1 port map( A => n3699, B => n3696, S => n677, Z => n3700);
   U4244 : MUX2_X1 port map( A => REGISTERS_21_4_port, B => REGISTERS_23_4_port
                           , S => n716, Z => n3701);
   U4245 : MUX2_X1 port map( A => REGISTERS_20_4_port, B => REGISTERS_22_4_port
                           , S => n716, Z => n3702);
   U4246 : MUX2_X1 port map( A => n3702, B => n3701, S => n750, Z => n3703);
   U4247 : MUX2_X1 port map( A => REGISTERS_17_4_port, B => REGISTERS_19_4_port
                           , S => n716, Z => n3704);
   U4248 : MUX2_X1 port map( A => REGISTERS_16_4_port, B => REGISTERS_18_4_port
                           , S => n716, Z => n3705);
   U4249 : MUX2_X1 port map( A => n3705, B => n3704, S => n750, Z => n3706);
   U4250 : MUX2_X1 port map( A => n3706, B => n3703, S => n677, Z => n3707);
   U4251 : MUX2_X1 port map( A => n3707, B => n3700, S => r3007_A_3_port, Z => 
                           n3708);
   U4252 : MUX2_X1 port map( A => REGISTERS_13_4_port, B => REGISTERS_15_4_port
                           , S => n716, Z => n3709);
   U4253 : MUX2_X1 port map( A => REGISTERS_12_4_port, B => REGISTERS_14_4_port
                           , S => n716, Z => n3710);
   U4254 : MUX2_X1 port map( A => n3710, B => n3709, S => n750, Z => n3711);
   U4255 : MUX2_X1 port map( A => REGISTERS_9_4_port, B => REGISTERS_11_4_port,
                           S => n716, Z => n3712);
   U4256 : MUX2_X1 port map( A => REGISTERS_8_4_port, B => REGISTERS_10_4_port,
                           S => n716, Z => n3713);
   U4257 : MUX2_X1 port map( A => n3713, B => n3712, S => n750, Z => n3714);
   U4258 : MUX2_X1 port map( A => n3714, B => n3711, S => n677, Z => n3715);
   U4259 : MUX2_X1 port map( A => REGISTERS_5_4_port, B => REGISTERS_7_4_port, 
                           S => n716, Z => n3716);
   U4260 : MUX2_X1 port map( A => REGISTERS_4_4_port, B => REGISTERS_6_4_port, 
                           S => n716, Z => n3717);
   U4261 : MUX2_X1 port map( A => n3717, B => n3716, S => n750, Z => n3718);
   U4262 : MUX2_X1 port map( A => REGISTERS_1_4_port, B => REGISTERS_3_4_port, 
                           S => n716, Z => n3719);
   U4263 : MUX2_X1 port map( A => REGISTERS_0_4_port, B => REGISTERS_2_4_port, 
                           S => n716, Z => n3720);
   U4264 : MUX2_X1 port map( A => n3720, B => n3719, S => n750, Z => n3721);
   U4265 : MUX2_X1 port map( A => n3721, B => n3718, S => n677, Z => n3722);
   U4266 : MUX2_X1 port map( A => n3722, B => n3715, S => r3007_A_3_port, Z => 
                           n3723);
   U4267 : MUX2_X1 port map( A => n3723, B => n3708, S => r3007_A_4_port, Z => 
                           n3724);
   U4268 : MUX2_X1 port map( A => n3724, B => n3693, S => ADD_RD1_5_port, Z => 
                           N4416);
   U4269 : MUX2_X1 port map( A => REGISTERS_37_5_port, B => REGISTERS_39_5_port
                           , S => n716, Z => n3725);
   U4270 : MUX2_X1 port map( A => REGISTERS_36_5_port, B => REGISTERS_38_5_port
                           , S => n716, Z => n3726);
   U4271 : MUX2_X1 port map( A => n3726, B => n3725, S => n750, Z => n3727);
   U4272 : MUX2_X1 port map( A => REGISTERS_33_5_port, B => REGISTERS_35_5_port
                           , S => n715, Z => n3728);
   U4273 : MUX2_X1 port map( A => REGISTERS_32_5_port, B => REGISTERS_34_5_port
                           , S => n715, Z => n3729);
   U4274 : MUX2_X1 port map( A => n3729, B => n3728, S => n750, Z => n3730);
   U4275 : MUX2_X1 port map( A => n3730, B => n3727, S => n677, Z => n3731);
   U4276 : MUX2_X1 port map( A => REGISTERS_29_5_port, B => REGISTERS_31_5_port
                           , S => n715, Z => n3732);
   U4277 : MUX2_X1 port map( A => REGISTERS_28_5_port, B => REGISTERS_30_5_port
                           , S => n715, Z => n3733);
   U4278 : MUX2_X1 port map( A => n3733, B => n3732, S => n749, Z => n3734);
   U4279 : MUX2_X1 port map( A => REGISTERS_25_5_port, B => REGISTERS_27_5_port
                           , S => n715, Z => n3735);
   U4280 : MUX2_X1 port map( A => REGISTERS_24_5_port, B => REGISTERS_26_5_port
                           , S => n715, Z => n3736);
   U4281 : MUX2_X1 port map( A => n3736, B => n3735, S => n749, Z => n3737);
   U4282 : MUX2_X1 port map( A => n3737, B => n3734, S => n677, Z => n3738);
   U4283 : MUX2_X1 port map( A => REGISTERS_21_5_port, B => REGISTERS_23_5_port
                           , S => n715, Z => n3739);
   U4284 : MUX2_X1 port map( A => REGISTERS_20_5_port, B => REGISTERS_22_5_port
                           , S => n715, Z => n3740);
   U4285 : MUX2_X1 port map( A => n3740, B => n3739, S => n749, Z => n3741);
   U4286 : MUX2_X1 port map( A => REGISTERS_17_5_port, B => REGISTERS_19_5_port
                           , S => n715, Z => n3742);
   U4287 : MUX2_X1 port map( A => REGISTERS_16_5_port, B => REGISTERS_18_5_port
                           , S => n715, Z => n3743);
   U4288 : MUX2_X1 port map( A => n3743, B => n3742, S => n749, Z => n3744);
   U4289 : MUX2_X1 port map( A => n3744, B => n3741, S => n677, Z => n3745);
   U4290 : MUX2_X1 port map( A => n3745, B => n3738, S => r3007_A_3_port, Z => 
                           n3746);
   U4291 : MUX2_X1 port map( A => REGISTERS_13_5_port, B => REGISTERS_15_5_port
                           , S => n715, Z => n3747);
   U4292 : MUX2_X1 port map( A => REGISTERS_12_5_port, B => REGISTERS_14_5_port
                           , S => n715, Z => n3748);
   U4293 : MUX2_X1 port map( A => n3748, B => n3747, S => n749, Z => n3749);
   U4294 : MUX2_X1 port map( A => REGISTERS_9_5_port, B => REGISTERS_11_5_port,
                           S => n715, Z => n3750);
   U4295 : MUX2_X1 port map( A => REGISTERS_8_5_port, B => REGISTERS_10_5_port,
                           S => n715, Z => n3751);
   U4296 : MUX2_X1 port map( A => n3751, B => n3750, S => n749, Z => n3752);
   U4297 : MUX2_X1 port map( A => n3752, B => n3749, S => n677, Z => n3753);
   U4298 : MUX2_X1 port map( A => REGISTERS_5_5_port, B => REGISTERS_7_5_port, 
                           S => n715, Z => n3754);
   U4299 : MUX2_X1 port map( A => REGISTERS_4_5_port, B => REGISTERS_6_5_port, 
                           S => n714, Z => n3755);
   U4300 : MUX2_X1 port map( A => n3755, B => n3754, S => n749, Z => n3756);
   U4301 : MUX2_X1 port map( A => REGISTERS_1_5_port, B => REGISTERS_3_5_port, 
                           S => n714, Z => n3757);
   U4302 : MUX2_X1 port map( A => REGISTERS_0_5_port, B => REGISTERS_2_5_port, 
                           S => n714, Z => n3758);
   U4303 : MUX2_X1 port map( A => n3758, B => n3757, S => n749, Z => n3759);
   U4304 : MUX2_X1 port map( A => n3759, B => n3756, S => n677, Z => n3760);
   U4305 : MUX2_X1 port map( A => n3760, B => n3753, S => r3007_A_3_port, Z => 
                           n3761);
   U4306 : MUX2_X1 port map( A => n3761, B => n3746, S => r3007_A_4_port, Z => 
                           n3762);
   U4307 : MUX2_X1 port map( A => n3762, B => n3731, S => ADD_RD1_5_port, Z => 
                           N4415);
   U4308 : MUX2_X1 port map( A => REGISTERS_37_6_port, B => REGISTERS_39_6_port
                           , S => n714, Z => n3763);
   U4309 : MUX2_X1 port map( A => REGISTERS_36_6_port, B => REGISTERS_38_6_port
                           , S => n714, Z => n3764);
   U4310 : MUX2_X1 port map( A => n3764, B => n3763, S => n749, Z => n3765);
   U4311 : MUX2_X1 port map( A => REGISTERS_33_6_port, B => REGISTERS_35_6_port
                           , S => n714, Z => n3766);
   U4312 : MUX2_X1 port map( A => REGISTERS_32_6_port, B => REGISTERS_34_6_port
                           , S => n714, Z => n3767);
   U4313 : MUX2_X1 port map( A => n3767, B => n3766, S => n749, Z => n3768);
   U4314 : MUX2_X1 port map( A => n3768, B => n3765, S => n677, Z => n3769);
   U4315 : MUX2_X1 port map( A => REGISTERS_29_6_port, B => REGISTERS_31_6_port
                           , S => n714, Z => n3770);
   U4316 : MUX2_X1 port map( A => REGISTERS_28_6_port, B => REGISTERS_30_6_port
                           , S => n714, Z => n3771);
   U4317 : MUX2_X1 port map( A => n3771, B => n3770, S => n749, Z => n3772);
   U4318 : MUX2_X1 port map( A => REGISTERS_25_6_port, B => REGISTERS_27_6_port
                           , S => n714, Z => n3773);
   U4319 : MUX2_X1 port map( A => REGISTERS_24_6_port, B => REGISTERS_26_6_port
                           , S => n714, Z => n3774);
   U4320 : MUX2_X1 port map( A => n3774, B => n3773, S => n749, Z => n3775);
   U4321 : MUX2_X1 port map( A => n3775, B => n3772, S => n677, Z => n3776);
   U4322 : MUX2_X1 port map( A => REGISTERS_21_6_port, B => REGISTERS_23_6_port
                           , S => n714, Z => n3777);
   U4323 : MUX2_X1 port map( A => REGISTERS_20_6_port, B => REGISTERS_22_6_port
                           , S => n714, Z => n3778);
   U4324 : MUX2_X1 port map( A => n3778, B => n3777, S => n749, Z => n3779);
   U4325 : MUX2_X1 port map( A => REGISTERS_17_6_port, B => REGISTERS_19_6_port
                           , S => n714, Z => n3780);
   U4326 : MUX2_X1 port map( A => REGISTERS_16_6_port, B => REGISTERS_18_6_port
                           , S => n714, Z => n3781);
   U4327 : MUX2_X1 port map( A => n3781, B => n3780, S => n749, Z => n3782);
   U4328 : MUX2_X1 port map( A => n3782, B => n3779, S => n677, Z => n3783);
   U4329 : MUX2_X1 port map( A => n3783, B => n3776, S => r3007_A_3_port, Z => 
                           n3784);
   U4330 : MUX2_X1 port map( A => REGISTERS_13_6_port, B => REGISTERS_15_6_port
                           , S => n713, Z => n3785);
   U4331 : MUX2_X1 port map( A => REGISTERS_12_6_port, B => REGISTERS_14_6_port
                           , S => n713, Z => n3786);
   U4332 : MUX2_X1 port map( A => n3786, B => n3785, S => n749, Z => n3787);
   U4333 : MUX2_X1 port map( A => REGISTERS_9_6_port, B => REGISTERS_11_6_port,
                           S => n713, Z => n3788);
   U4334 : MUX2_X1 port map( A => REGISTERS_8_6_port, B => REGISTERS_10_6_port,
                           S => n713, Z => n3789);
   U4335 : MUX2_X1 port map( A => n3789, B => n3788, S => n748, Z => n3790);
   U4336 : MUX2_X1 port map( A => n3790, B => n3787, S => n677, Z => n3791);
   U4337 : MUX2_X1 port map( A => REGISTERS_5_6_port, B => REGISTERS_7_6_port, 
                           S => n713, Z => n3792);
   U4338 : MUX2_X1 port map( A => REGISTERS_4_6_port, B => REGISTERS_6_6_port, 
                           S => n713, Z => n3793);
   U4339 : MUX2_X1 port map( A => n3793, B => n3792, S => n748, Z => n3794);
   U4340 : MUX2_X1 port map( A => REGISTERS_1_6_port, B => REGISTERS_3_6_port, 
                           S => n713, Z => n3795);
   U4341 : MUX2_X1 port map( A => REGISTERS_0_6_port, B => REGISTERS_2_6_port, 
                           S => n713, Z => n3796);
   U4342 : MUX2_X1 port map( A => n3796, B => n3795, S => n748, Z => n3797);
   U4343 : MUX2_X1 port map( A => n3797, B => n3794, S => n677, Z => n3798);
   U4344 : MUX2_X1 port map( A => n3798, B => n3791, S => r3007_A_3_port, Z => 
                           n3799);
   U4345 : MUX2_X1 port map( A => n3799, B => n3784, S => r3007_A_4_port, Z => 
                           n3800);
   U4346 : MUX2_X1 port map( A => n3800, B => n3769, S => ADD_RD1_5_port, Z => 
                           N4414);
   U4347 : MUX2_X1 port map( A => REGISTERS_37_7_port, B => REGISTERS_39_7_port
                           , S => n713, Z => n3801);
   U4348 : MUX2_X1 port map( A => REGISTERS_36_7_port, B => REGISTERS_38_7_port
                           , S => n713, Z => n3802);
   U4349 : MUX2_X1 port map( A => n3802, B => n3801, S => n748, Z => n3803);
   U4350 : MUX2_X1 port map( A => REGISTERS_33_7_port, B => REGISTERS_35_7_port
                           , S => n713, Z => n3804);
   U4351 : MUX2_X1 port map( A => REGISTERS_32_7_port, B => REGISTERS_34_7_port
                           , S => n713, Z => n3805);
   U4352 : MUX2_X1 port map( A => n3805, B => n3804, S => n748, Z => n3806);
   U4353 : MUX2_X1 port map( A => n3806, B => n3803, S => n676, Z => n3807);
   U4354 : MUX2_X1 port map( A => REGISTERS_29_7_port, B => REGISTERS_31_7_port
                           , S => n713, Z => n3808);
   U4355 : MUX2_X1 port map( A => REGISTERS_28_7_port, B => REGISTERS_30_7_port
                           , S => n713, Z => n3809);
   U4356 : MUX2_X1 port map( A => n3809, B => n3808, S => n748, Z => n3810);
   U4357 : MUX2_X1 port map( A => REGISTERS_25_7_port, B => REGISTERS_27_7_port
                           , S => n713, Z => n3811);
   U4358 : MUX2_X1 port map( A => REGISTERS_24_7_port, B => REGISTERS_26_7_port
                           , S => n712, Z => n3812);
   U4359 : MUX2_X1 port map( A => n3812, B => n3811, S => n748, Z => n3813);
   U4360 : MUX2_X1 port map( A => n3813, B => n3810, S => n676, Z => n3814);
   U4361 : MUX2_X1 port map( A => REGISTERS_21_7_port, B => REGISTERS_23_7_port
                           , S => n712, Z => n3815);
   U4362 : MUX2_X1 port map( A => REGISTERS_20_7_port, B => REGISTERS_22_7_port
                           , S => n712, Z => n3816);
   U4363 : MUX2_X1 port map( A => n3816, B => n3815, S => n748, Z => n3817);
   U4364 : MUX2_X1 port map( A => REGISTERS_17_7_port, B => REGISTERS_19_7_port
                           , S => n712, Z => n3818);
   U4365 : MUX2_X1 port map( A => REGISTERS_16_7_port, B => REGISTERS_18_7_port
                           , S => n712, Z => n3819);
   U4366 : MUX2_X1 port map( A => n3819, B => n3818, S => n748, Z => n3820);
   U4367 : MUX2_X1 port map( A => n3820, B => n3817, S => n676, Z => n3821);
   U4368 : MUX2_X1 port map( A => n3821, B => n3814, S => r3007_A_3_port, Z => 
                           n3822);
   U4369 : MUX2_X1 port map( A => REGISTERS_13_7_port, B => REGISTERS_15_7_port
                           , S => n712, Z => n3823);
   U4370 : MUX2_X1 port map( A => REGISTERS_12_7_port, B => REGISTERS_14_7_port
                           , S => n712, Z => n3824);
   U4371 : MUX2_X1 port map( A => n3824, B => n3823, S => n748, Z => n3825);
   U4372 : MUX2_X1 port map( A => REGISTERS_9_7_port, B => REGISTERS_11_7_port,
                           S => n712, Z => n3826);
   U4373 : MUX2_X1 port map( A => REGISTERS_8_7_port, B => REGISTERS_10_7_port,
                           S => n712, Z => n3827);
   U4374 : MUX2_X1 port map( A => n3827, B => n3826, S => n748, Z => n3828);
   U4375 : MUX2_X1 port map( A => n3828, B => n3825, S => n676, Z => n3829);
   U4376 : MUX2_X1 port map( A => REGISTERS_5_7_port, B => REGISTERS_7_7_port, 
                           S => n712, Z => n3830);
   U4377 : MUX2_X1 port map( A => REGISTERS_4_7_port, B => REGISTERS_6_7_port, 
                           S => n712, Z => n3831);
   U4378 : MUX2_X1 port map( A => n3831, B => n3830, S => n748, Z => n3832);
   U4379 : MUX2_X1 port map( A => REGISTERS_1_7_port, B => REGISTERS_3_7_port, 
                           S => n712, Z => n3833);
   U4380 : MUX2_X1 port map( A => REGISTERS_0_7_port, B => REGISTERS_2_7_port, 
                           S => n712, Z => n3834);
   U4381 : MUX2_X1 port map( A => n3834, B => n3833, S => n748, Z => n3835);
   U4382 : MUX2_X1 port map( A => n3835, B => n3832, S => n676, Z => n3836);
   U4383 : MUX2_X1 port map( A => n3836, B => n3829, S => r3007_A_3_port, Z => 
                           n3837);
   U4384 : MUX2_X1 port map( A => n3837, B => n3822, S => r3007_A_4_port, Z => 
                           n3838);
   U4385 : MUX2_X1 port map( A => n3838, B => n3807, S => ADD_RD1_5_port, Z => 
                           N4413);
   U4386 : MUX2_X1 port map( A => REGISTERS_37_8_port, B => REGISTERS_39_8_port
                           , S => n712, Z => n3839);
   U4387 : MUX2_X1 port map( A => REGISTERS_36_8_port, B => REGISTERS_38_8_port
                           , S => n712, Z => n3840);
   U4388 : MUX2_X1 port map( A => n3840, B => n3839, S => n748, Z => n3841);
   U4389 : MUX2_X1 port map( A => REGISTERS_33_8_port, B => REGISTERS_35_8_port
                           , S => n711, Z => n3842);
   U4390 : MUX2_X1 port map( A => REGISTERS_32_8_port, B => REGISTERS_34_8_port
                           , S => n711, Z => n3843);
   U4391 : MUX2_X1 port map( A => n3843, B => n3842, S => n748, Z => n3844);
   U4392 : MUX2_X1 port map( A => n3844, B => n3841, S => n676, Z => n3845);
   U4393 : MUX2_X1 port map( A => REGISTERS_29_8_port, B => REGISTERS_31_8_port
                           , S => n711, Z => n3846);
   U4394 : MUX2_X1 port map( A => REGISTERS_28_8_port, B => REGISTERS_30_8_port
                           , S => n711, Z => n3847);
   U4395 : MUX2_X1 port map( A => n3847, B => n3846, S => n747, Z => n3848);
   U4396 : MUX2_X1 port map( A => REGISTERS_25_8_port, B => REGISTERS_27_8_port
                           , S => n711, Z => n3849);
   U4397 : MUX2_X1 port map( A => REGISTERS_24_8_port, B => REGISTERS_26_8_port
                           , S => n711, Z => n3850);
   U4398 : MUX2_X1 port map( A => n3850, B => n3849, S => n747, Z => n3851);
   U4399 : MUX2_X1 port map( A => n3851, B => n3848, S => n676, Z => n3852);
   U4400 : MUX2_X1 port map( A => REGISTERS_21_8_port, B => REGISTERS_23_8_port
                           , S => n711, Z => n3853);
   U4401 : MUX2_X1 port map( A => REGISTERS_20_8_port, B => REGISTERS_22_8_port
                           , S => n711, Z => n3854);
   U4402 : MUX2_X1 port map( A => n3854, B => n3853, S => n747, Z => n3855);
   U4403 : MUX2_X1 port map( A => REGISTERS_17_8_port, B => REGISTERS_19_8_port
                           , S => n711, Z => n3856);
   U4404 : MUX2_X1 port map( A => REGISTERS_16_8_port, B => REGISTERS_18_8_port
                           , S => n711, Z => n3857);
   U4405 : MUX2_X1 port map( A => n3857, B => n3856, S => n747, Z => n3858);
   U4406 : MUX2_X1 port map( A => n3858, B => n3855, S => n676, Z => n3859);
   U4407 : MUX2_X1 port map( A => n3859, B => n3852, S => r3007_A_3_port, Z => 
                           n3860);
   U4408 : MUX2_X1 port map( A => REGISTERS_13_8_port, B => REGISTERS_15_8_port
                           , S => n711, Z => n3861);
   U4409 : MUX2_X1 port map( A => REGISTERS_12_8_port, B => REGISTERS_14_8_port
                           , S => n711, Z => n3862);
   U4410 : MUX2_X1 port map( A => n3862, B => n3861, S => n747, Z => n3863);
   U4411 : MUX2_X1 port map( A => REGISTERS_9_8_port, B => REGISTERS_11_8_port,
                           S => n711, Z => n3864);
   U4412 : MUX2_X1 port map( A => REGISTERS_8_8_port, B => REGISTERS_10_8_port,
                           S => n711, Z => n3865);
   U4413 : MUX2_X1 port map( A => n3865, B => n3864, S => n747, Z => n3866);
   U4414 : MUX2_X1 port map( A => n3866, B => n3863, S => n676, Z => n3867);
   U4415 : MUX2_X1 port map( A => REGISTERS_5_8_port, B => REGISTERS_7_8_port, 
                           S => n711, Z => n3868);
   U4416 : MUX2_X1 port map( A => REGISTERS_4_8_port, B => REGISTERS_6_8_port, 
                           S => n710, Z => n3869);
   U4417 : MUX2_X1 port map( A => n3869, B => n3868, S => n747, Z => n3870);
   U4418 : MUX2_X1 port map( A => REGISTERS_1_8_port, B => REGISTERS_3_8_port, 
                           S => n710, Z => n3871);
   U4419 : MUX2_X1 port map( A => REGISTERS_0_8_port, B => REGISTERS_2_8_port, 
                           S => n710, Z => n3872);
   U4420 : MUX2_X1 port map( A => n3872, B => n3871, S => n747, Z => n3873);
   U4421 : MUX2_X1 port map( A => n3873, B => n3870, S => n676, Z => n3874);
   U4422 : MUX2_X1 port map( A => n3874, B => n3867, S => r3007_A_3_port, Z => 
                           n3875);
   U4423 : MUX2_X1 port map( A => n3875, B => n3860, S => r3007_A_4_port, Z => 
                           n3876);
   U4424 : MUX2_X1 port map( A => n3876, B => n3845, S => ADD_RD1_5_port, Z => 
                           N4412);
   U4425 : MUX2_X1 port map( A => REGISTERS_37_9_port, B => REGISTERS_39_9_port
                           , S => n710, Z => n3877);
   U4426 : MUX2_X1 port map( A => REGISTERS_36_9_port, B => REGISTERS_38_9_port
                           , S => n710, Z => n3878);
   U4427 : MUX2_X1 port map( A => n3878, B => n3877, S => n747, Z => n3879);
   U4428 : MUX2_X1 port map( A => REGISTERS_33_9_port, B => REGISTERS_35_9_port
                           , S => n710, Z => n3880);
   U4429 : MUX2_X1 port map( A => REGISTERS_32_9_port, B => REGISTERS_34_9_port
                           , S => n710, Z => n3881);
   U4430 : MUX2_X1 port map( A => n3881, B => n3880, S => n747, Z => n3882);
   U4431 : MUX2_X1 port map( A => n3882, B => n3879, S => n676, Z => n3883);
   U4432 : MUX2_X1 port map( A => REGISTERS_29_9_port, B => REGISTERS_31_9_port
                           , S => n710, Z => n3884);
   U4433 : MUX2_X1 port map( A => REGISTERS_28_9_port, B => REGISTERS_30_9_port
                           , S => n710, Z => n3885);
   U4434 : MUX2_X1 port map( A => n3885, B => n3884, S => n747, Z => n3886);
   U4435 : MUX2_X1 port map( A => REGISTERS_25_9_port, B => REGISTERS_27_9_port
                           , S => n710, Z => n3887);
   U4436 : MUX2_X1 port map( A => REGISTERS_24_9_port, B => REGISTERS_26_9_port
                           , S => n710, Z => n3888);
   U4437 : MUX2_X1 port map( A => n3888, B => n3887, S => n747, Z => n3889);
   U4438 : MUX2_X1 port map( A => n3889, B => n3886, S => n676, Z => n3890);
   U4439 : MUX2_X1 port map( A => REGISTERS_21_9_port, B => REGISTERS_23_9_port
                           , S => n710, Z => n3891);
   U4440 : MUX2_X1 port map( A => REGISTERS_20_9_port, B => REGISTERS_22_9_port
                           , S => n710, Z => n3892);
   U4441 : MUX2_X1 port map( A => n3892, B => n3891, S => n747, Z => n3893);
   U4442 : MUX2_X1 port map( A => REGISTERS_17_9_port, B => REGISTERS_19_9_port
                           , S => n710, Z => n3894);
   U4443 : MUX2_X1 port map( A => REGISTERS_16_9_port, B => REGISTERS_18_9_port
                           , S => n710, Z => n3895);
   U4444 : MUX2_X1 port map( A => n3895, B => n3894, S => n747, Z => n3896);
   U4445 : MUX2_X1 port map( A => n3896, B => n3893, S => n676, Z => n3897);
   U4446 : MUX2_X1 port map( A => n3897, B => n3890, S => r3007_A_3_port, Z => 
                           n3898);
   U4447 : MUX2_X1 port map( A => REGISTERS_13_9_port, B => REGISTERS_15_9_port
                           , S => n709, Z => n3899);
   U4448 : MUX2_X1 port map( A => REGISTERS_12_9_port, B => REGISTERS_14_9_port
                           , S => n709, Z => n3900);
   U4449 : MUX2_X1 port map( A => n3900, B => n3899, S => n747, Z => n3901);
   U4450 : MUX2_X1 port map( A => REGISTERS_9_9_port, B => REGISTERS_11_9_port,
                           S => n709, Z => n3902);
   U4451 : MUX2_X1 port map( A => REGISTERS_8_9_port, B => REGISTERS_10_9_port,
                           S => n709, Z => n3903);
   U4452 : MUX2_X1 port map( A => n3903, B => n3902, S => n746, Z => n3904);
   U4453 : MUX2_X1 port map( A => n3904, B => n3901, S => n676, Z => n3905);
   U4454 : MUX2_X1 port map( A => REGISTERS_5_9_port, B => REGISTERS_7_9_port, 
                           S => n709, Z => n3906);
   U4455 : MUX2_X1 port map( A => REGISTERS_4_9_port, B => REGISTERS_6_9_port, 
                           S => n709, Z => n3907);
   U4456 : MUX2_X1 port map( A => n3907, B => n3906, S => n746, Z => n3908);
   U4457 : MUX2_X1 port map( A => REGISTERS_1_9_port, B => REGISTERS_3_9_port, 
                           S => n709, Z => n3909);
   U4458 : MUX2_X1 port map( A => REGISTERS_0_9_port, B => REGISTERS_2_9_port, 
                           S => n709, Z => n3910);
   U4459 : MUX2_X1 port map( A => n3910, B => n3909, S => n746, Z => n3911);
   U4460 : MUX2_X1 port map( A => n3911, B => n3908, S => n675, Z => n3912);
   U4461 : MUX2_X1 port map( A => n3912, B => n3905, S => r3007_A_3_port, Z => 
                           n3913);
   U4462 : MUX2_X1 port map( A => n3913, B => n3898, S => r3007_A_4_port, Z => 
                           n3914);
   U4463 : MUX2_X1 port map( A => n3914, B => n3883, S => ADD_RD1_5_port, Z => 
                           N4411);
   U4464 : MUX2_X1 port map( A => REGISTERS_37_10_port, B => 
                           REGISTERS_39_10_port, S => n709, Z => n3915);
   U4465 : MUX2_X1 port map( A => REGISTERS_36_10_port, B => 
                           REGISTERS_38_10_port, S => n709, Z => n3916);
   U4466 : MUX2_X1 port map( A => n3916, B => n3915, S => n746, Z => n3917);
   U4467 : MUX2_X1 port map( A => REGISTERS_33_10_port, B => 
                           REGISTERS_35_10_port, S => n709, Z => n3918);
   U4468 : MUX2_X1 port map( A => REGISTERS_32_10_port, B => 
                           REGISTERS_34_10_port, S => n709, Z => n3919);
   U4469 : MUX2_X1 port map( A => n3919, B => n3918, S => n746, Z => n3920);
   U4470 : MUX2_X1 port map( A => n3920, B => n3917, S => n675, Z => n3921);
   U4471 : MUX2_X1 port map( A => REGISTERS_29_10_port, B => 
                           REGISTERS_31_10_port, S => n709, Z => n3922);
   U4472 : MUX2_X1 port map( A => REGISTERS_28_10_port, B => 
                           REGISTERS_30_10_port, S => n709, Z => n3923);
   U4473 : MUX2_X1 port map( A => n3923, B => n3922, S => n746, Z => n3924);
   U4474 : MUX2_X1 port map( A => REGISTERS_25_10_port, B => 
                           REGISTERS_27_10_port, S => n709, Z => n3925);
   U4475 : MUX2_X1 port map( A => REGISTERS_24_10_port, B => 
                           REGISTERS_26_10_port, S => n708, Z => n3926);
   U4476 : MUX2_X1 port map( A => n3926, B => n3925, S => n746, Z => n3927);
   U4477 : MUX2_X1 port map( A => n3927, B => n3924, S => n675, Z => n3928);
   U4478 : MUX2_X1 port map( A => REGISTERS_21_10_port, B => 
                           REGISTERS_23_10_port, S => n708, Z => n3929);
   U4479 : MUX2_X1 port map( A => REGISTERS_20_10_port, B => 
                           REGISTERS_22_10_port, S => n708, Z => n3930);
   U4480 : MUX2_X1 port map( A => n3930, B => n3929, S => n746, Z => n3931);
   U4481 : MUX2_X1 port map( A => REGISTERS_17_10_port, B => 
                           REGISTERS_19_10_port, S => n708, Z => n3932);
   U4482 : MUX2_X1 port map( A => REGISTERS_16_10_port, B => 
                           REGISTERS_18_10_port, S => n708, Z => n3933);
   U4483 : MUX2_X1 port map( A => n3933, B => n3932, S => n746, Z => n3934);
   U4484 : MUX2_X1 port map( A => n3934, B => n3931, S => n675, Z => n3935);
   U4485 : MUX2_X1 port map( A => n3935, B => n3928, S => r3007_A_3_port, Z => 
                           n3936);
   U4486 : MUX2_X1 port map( A => REGISTERS_13_10_port, B => 
                           REGISTERS_15_10_port, S => n708, Z => n3937);
   U4487 : MUX2_X1 port map( A => REGISTERS_12_10_port, B => 
                           REGISTERS_14_10_port, S => n708, Z => n3938);
   U4488 : MUX2_X1 port map( A => n3938, B => n3937, S => n746, Z => n3939);
   U4489 : MUX2_X1 port map( A => REGISTERS_9_10_port, B => 
                           REGISTERS_11_10_port, S => n708, Z => n3940);
   U4490 : MUX2_X1 port map( A => REGISTERS_8_10_port, B => 
                           REGISTERS_10_10_port, S => n708, Z => n3941);
   U4491 : MUX2_X1 port map( A => n3941, B => n3940, S => n746, Z => n3942);
   U4492 : MUX2_X1 port map( A => n3942, B => n3939, S => n675, Z => n3943);
   U4493 : MUX2_X1 port map( A => REGISTERS_5_10_port, B => REGISTERS_7_10_port
                           , S => n708, Z => n3944);
   U4494 : MUX2_X1 port map( A => REGISTERS_4_10_port, B => REGISTERS_6_10_port
                           , S => n708, Z => n3945);
   U4495 : MUX2_X1 port map( A => n3945, B => n3944, S => n746, Z => n3946);
   U4496 : MUX2_X1 port map( A => REGISTERS_1_10_port, B => REGISTERS_3_10_port
                           , S => n708, Z => n3947);
   U4497 : MUX2_X1 port map( A => REGISTERS_0_10_port, B => REGISTERS_2_10_port
                           , S => n708, Z => n3948);
   U4498 : MUX2_X1 port map( A => n3948, B => n3947, S => n746, Z => n3949);
   U4499 : MUX2_X1 port map( A => n3949, B => n3946, S => n675, Z => n3950);
   U4500 : MUX2_X1 port map( A => n3950, B => n3943, S => r3007_A_3_port, Z => 
                           n3951);
   U4501 : MUX2_X1 port map( A => n3951, B => n3936, S => r3007_A_4_port, Z => 
                           n3952);
   U4502 : MUX2_X1 port map( A => n3952, B => n3921, S => ADD_RD1_5_port, Z => 
                           N4410);
   U4503 : MUX2_X1 port map( A => REGISTERS_37_11_port, B => 
                           REGISTERS_39_11_port, S => n708, Z => n3953);
   U4504 : MUX2_X1 port map( A => REGISTERS_36_11_port, B => 
                           REGISTERS_38_11_port, S => n708, Z => n3954);
   U4505 : MUX2_X1 port map( A => n3954, B => n3953, S => n746, Z => n3955);
   U4506 : MUX2_X1 port map( A => REGISTERS_33_11_port, B => 
                           REGISTERS_35_11_port, S => n707, Z => n3956);
   U4507 : MUX2_X1 port map( A => REGISTERS_32_11_port, B => 
                           REGISTERS_34_11_port, S => n707, Z => n3957);
   U4508 : MUX2_X1 port map( A => n3957, B => n3956, S => n746, Z => n3958);
   U4509 : MUX2_X1 port map( A => n3958, B => n3955, S => n675, Z => n3959);
   U4510 : MUX2_X1 port map( A => REGISTERS_29_11_port, B => 
                           REGISTERS_31_11_port, S => n707, Z => n3960);
   U4511 : MUX2_X1 port map( A => REGISTERS_28_11_port, B => 
                           REGISTERS_30_11_port, S => n707, Z => n3961);
   U4512 : MUX2_X1 port map( A => n3961, B => n3960, S => n745, Z => n3962);
   U4513 : MUX2_X1 port map( A => REGISTERS_25_11_port, B => 
                           REGISTERS_27_11_port, S => n707, Z => n3963);
   U4514 : MUX2_X1 port map( A => REGISTERS_24_11_port, B => 
                           REGISTERS_26_11_port, S => n707, Z => n3964);
   U4515 : MUX2_X1 port map( A => n3964, B => n3963, S => n745, Z => n3965);
   U4516 : MUX2_X1 port map( A => n3965, B => n3962, S => n675, Z => n3966);
   U4517 : MUX2_X1 port map( A => REGISTERS_21_11_port, B => 
                           REGISTERS_23_11_port, S => n707, Z => n3967);
   U4518 : MUX2_X1 port map( A => REGISTERS_20_11_port, B => 
                           REGISTERS_22_11_port, S => n707, Z => n3968);
   U4519 : MUX2_X1 port map( A => n3968, B => n3967, S => n745, Z => n3969);
   U4520 : MUX2_X1 port map( A => REGISTERS_17_11_port, B => 
                           REGISTERS_19_11_port, S => n707, Z => n3970);
   U4521 : MUX2_X1 port map( A => REGISTERS_16_11_port, B => 
                           REGISTERS_18_11_port, S => n707, Z => n3971);
   U4522 : MUX2_X1 port map( A => n3971, B => n3970, S => n745, Z => n3972);
   U4523 : MUX2_X1 port map( A => n3972, B => n3969, S => n675, Z => n3973);
   U4524 : MUX2_X1 port map( A => n3973, B => n3966, S => r3007_A_3_port, Z => 
                           n3974);
   U4525 : MUX2_X1 port map( A => REGISTERS_13_11_port, B => 
                           REGISTERS_15_11_port, S => n707, Z => n3975);
   U4526 : MUX2_X1 port map( A => REGISTERS_12_11_port, B => 
                           REGISTERS_14_11_port, S => n707, Z => n3976);
   U4527 : MUX2_X1 port map( A => n3976, B => n3975, S => n745, Z => n3977);
   U4528 : MUX2_X1 port map( A => REGISTERS_9_11_port, B => 
                           REGISTERS_11_11_port, S => n707, Z => n3978);
   U4529 : MUX2_X1 port map( A => REGISTERS_8_11_port, B => 
                           REGISTERS_10_11_port, S => n707, Z => n3979);
   U4530 : MUX2_X1 port map( A => n3979, B => n3978, S => n745, Z => n3980);
   U4531 : MUX2_X1 port map( A => n3980, B => n3977, S => n675, Z => n3981);
   U4532 : MUX2_X1 port map( A => REGISTERS_5_11_port, B => REGISTERS_7_11_port
                           , S => n707, Z => n3982);
   U4533 : MUX2_X1 port map( A => REGISTERS_4_11_port, B => REGISTERS_6_11_port
                           , S => n706, Z => n3983);
   U4534 : MUX2_X1 port map( A => n3983, B => n3982, S => n745, Z => n3984);
   U4535 : MUX2_X1 port map( A => REGISTERS_1_11_port, B => REGISTERS_3_11_port
                           , S => n706, Z => n3985);
   U4536 : MUX2_X1 port map( A => REGISTERS_0_11_port, B => REGISTERS_2_11_port
                           , S => n706, Z => n3986);
   U4537 : MUX2_X1 port map( A => n3986, B => n3985, S => n745, Z => n3987);
   U4538 : MUX2_X1 port map( A => n3987, B => n3984, S => n675, Z => n3988);
   U4539 : MUX2_X1 port map( A => n3988, B => n3981, S => r3007_A_3_port, Z => 
                           n3989);
   U4540 : MUX2_X1 port map( A => n3989, B => n3974, S => r3007_A_4_port, Z => 
                           n3990);
   U4541 : MUX2_X1 port map( A => n3990, B => n3959, S => ADD_RD1_5_port, Z => 
                           N4409);
   U4542 : MUX2_X1 port map( A => REGISTERS_37_12_port, B => 
                           REGISTERS_39_12_port, S => n706, Z => n3991);
   U4543 : MUX2_X1 port map( A => REGISTERS_36_12_port, B => 
                           REGISTERS_38_12_port, S => n706, Z => n3992);
   U4544 : MUX2_X1 port map( A => n3992, B => n3991, S => n745, Z => n3993);
   U4545 : MUX2_X1 port map( A => REGISTERS_33_12_port, B => 
                           REGISTERS_35_12_port, S => n706, Z => n3994);
   U4546 : MUX2_X1 port map( A => REGISTERS_32_12_port, B => 
                           REGISTERS_34_12_port, S => n706, Z => n3995);
   U4547 : MUX2_X1 port map( A => n3995, B => n3994, S => n745, Z => n3996);
   U4548 : MUX2_X1 port map( A => n3996, B => n3993, S => n675, Z => n3997);
   U4549 : MUX2_X1 port map( A => REGISTERS_29_12_port, B => 
                           REGISTERS_31_12_port, S => n706, Z => n3998);
   U4550 : MUX2_X1 port map( A => REGISTERS_28_12_port, B => 
                           REGISTERS_30_12_port, S => n706, Z => n3999);
   U4551 : MUX2_X1 port map( A => n3999, B => n3998, S => n745, Z => n4000);
   U4552 : MUX2_X1 port map( A => REGISTERS_25_12_port, B => 
                           REGISTERS_27_12_port, S => n706, Z => n4001);
   U4553 : MUX2_X1 port map( A => REGISTERS_24_12_port, B => 
                           REGISTERS_26_12_port, S => n706, Z => n4002);
   U4554 : MUX2_X1 port map( A => n4002, B => n4001, S => n745, Z => n4003);
   U4555 : MUX2_X1 port map( A => n4003, B => n4000, S => n675, Z => n4004);
   U4556 : MUX2_X1 port map( A => REGISTERS_21_12_port, B => 
                           REGISTERS_23_12_port, S => n706, Z => n4005);
   U4557 : MUX2_X1 port map( A => REGISTERS_20_12_port, B => 
                           REGISTERS_22_12_port, S => n706, Z => n4006);
   U4558 : MUX2_X1 port map( A => n4006, B => n4005, S => n745, Z => n4007);
   U4559 : MUX2_X1 port map( A => REGISTERS_17_12_port, B => 
                           REGISTERS_19_12_port, S => n706, Z => n4008);
   U4560 : MUX2_X1 port map( A => REGISTERS_16_12_port, B => 
                           REGISTERS_18_12_port, S => n706, Z => n4009);
   U4561 : MUX2_X1 port map( A => n4009, B => n4008, S => n745, Z => n4010);
   U4562 : MUX2_X1 port map( A => n4010, B => n4007, S => n675, Z => n4011);
   U4563 : MUX2_X1 port map( A => n4011, B => n4004, S => r3007_A_3_port, Z => 
                           n4012);
   U4564 : MUX2_X1 port map( A => REGISTERS_13_12_port, B => 
                           REGISTERS_15_12_port, S => n705, Z => n4013);
   U4565 : MUX2_X1 port map( A => REGISTERS_12_12_port, B => 
                           REGISTERS_14_12_port, S => n705, Z => n4014);
   U4566 : MUX2_X1 port map( A => n4014, B => n4013, S => n745, Z => n4015);
   U4567 : MUX2_X1 port map( A => REGISTERS_9_12_port, B => 
                           REGISTERS_11_12_port, S => n705, Z => n4016);
   U4568 : MUX2_X1 port map( A => REGISTERS_8_12_port, B => 
                           REGISTERS_10_12_port, S => n705, Z => n4017);
   U4569 : MUX2_X1 port map( A => n4017, B => n4016, S => n744, Z => n4018);
   U4570 : MUX2_X1 port map( A => n4018, B => n4015, S => n674, Z => n4019);
   U4571 : MUX2_X1 port map( A => REGISTERS_5_12_port, B => REGISTERS_7_12_port
                           , S => n705, Z => n4020);
   U4572 : MUX2_X1 port map( A => REGISTERS_4_12_port, B => REGISTERS_6_12_port
                           , S => n705, Z => n4021);
   U4573 : MUX2_X1 port map( A => n4021, B => n4020, S => n744, Z => n4022);
   U4574 : MUX2_X1 port map( A => REGISTERS_1_12_port, B => REGISTERS_3_12_port
                           , S => n705, Z => n4023);
   U4575 : MUX2_X1 port map( A => REGISTERS_0_12_port, B => REGISTERS_2_12_port
                           , S => n705, Z => n4024);
   U4576 : MUX2_X1 port map( A => n4024, B => n4023, S => n744, Z => n4025);
   U4577 : MUX2_X1 port map( A => n4025, B => n4022, S => n674, Z => n4026);
   U4578 : MUX2_X1 port map( A => n4026, B => n4019, S => r3007_A_3_port, Z => 
                           n4027);
   U4579 : MUX2_X1 port map( A => n4027, B => n4012, S => r3007_A_4_port, Z => 
                           n4028);
   U4580 : MUX2_X1 port map( A => n4028, B => n3997, S => ADD_RD1_5_port, Z => 
                           N4408);
   U4581 : MUX2_X1 port map( A => REGISTERS_37_13_port, B => 
                           REGISTERS_39_13_port, S => n705, Z => n4029);
   U4582 : MUX2_X1 port map( A => REGISTERS_36_13_port, B => 
                           REGISTERS_38_13_port, S => n705, Z => n4030);
   U4583 : MUX2_X1 port map( A => n4030, B => n4029, S => n744, Z => n4031);
   U4584 : MUX2_X1 port map( A => REGISTERS_33_13_port, B => 
                           REGISTERS_35_13_port, S => n705, Z => n4032);
   U4585 : MUX2_X1 port map( A => REGISTERS_32_13_port, B => 
                           REGISTERS_34_13_port, S => n705, Z => n4033);
   U4586 : MUX2_X1 port map( A => n4033, B => n4032, S => n744, Z => n4034);
   U4587 : MUX2_X1 port map( A => n4034, B => n4031, S => n674, Z => n4035);
   U4588 : MUX2_X1 port map( A => REGISTERS_29_13_port, B => 
                           REGISTERS_31_13_port, S => n705, Z => n4036);
   U4589 : MUX2_X1 port map( A => REGISTERS_28_13_port, B => 
                           REGISTERS_30_13_port, S => n705, Z => n4037);
   U4590 : MUX2_X1 port map( A => n4037, B => n4036, S => n744, Z => n4038);
   U4591 : MUX2_X1 port map( A => REGISTERS_25_13_port, B => 
                           REGISTERS_27_13_port, S => n705, Z => n4039);
   U4592 : MUX2_X1 port map( A => REGISTERS_24_13_port, B => 
                           REGISTERS_26_13_port, S => n704, Z => n4040);
   U4593 : MUX2_X1 port map( A => n4040, B => n4039, S => n744, Z => n4041);
   U4594 : MUX2_X1 port map( A => n4041, B => n4038, S => n674, Z => n4042);
   U4595 : MUX2_X1 port map( A => REGISTERS_21_13_port, B => 
                           REGISTERS_23_13_port, S => n704, Z => n4043);
   U4596 : MUX2_X1 port map( A => REGISTERS_20_13_port, B => 
                           REGISTERS_22_13_port, S => n704, Z => n4044);
   U4597 : MUX2_X1 port map( A => n4044, B => n4043, S => n744, Z => n4045);
   U4598 : MUX2_X1 port map( A => REGISTERS_17_13_port, B => 
                           REGISTERS_19_13_port, S => n704, Z => n4046);
   U4599 : MUX2_X1 port map( A => REGISTERS_16_13_port, B => 
                           REGISTERS_18_13_port, S => n704, Z => n4047);
   U4600 : MUX2_X1 port map( A => n4047, B => n4046, S => n744, Z => n4048);
   U4601 : MUX2_X1 port map( A => n4048, B => n4045, S => n674, Z => n4049);
   U4602 : MUX2_X1 port map( A => n4049, B => n4042, S => r3007_A_3_port, Z => 
                           n4050);
   U4603 : MUX2_X1 port map( A => REGISTERS_13_13_port, B => 
                           REGISTERS_15_13_port, S => n704, Z => n4051);
   U4604 : MUX2_X1 port map( A => REGISTERS_12_13_port, B => 
                           REGISTERS_14_13_port, S => n704, Z => n4052);
   U4605 : MUX2_X1 port map( A => n4052, B => n4051, S => n744, Z => n4053);
   U4606 : MUX2_X1 port map( A => REGISTERS_9_13_port, B => 
                           REGISTERS_11_13_port, S => n704, Z => n4054);
   U4607 : MUX2_X1 port map( A => REGISTERS_8_13_port, B => 
                           REGISTERS_10_13_port, S => n704, Z => n4055);
   U4608 : MUX2_X1 port map( A => n4055, B => n4054, S => n744, Z => n4056);
   U4609 : MUX2_X1 port map( A => n4056, B => n4053, S => n674, Z => n4057);
   U4610 : MUX2_X1 port map( A => REGISTERS_5_13_port, B => REGISTERS_7_13_port
                           , S => n704, Z => n4058);
   U4611 : MUX2_X1 port map( A => REGISTERS_4_13_port, B => REGISTERS_6_13_port
                           , S => n704, Z => n4059);
   U4612 : MUX2_X1 port map( A => n4059, B => n4058, S => n744, Z => n4060);
   U4613 : MUX2_X1 port map( A => REGISTERS_1_13_port, B => REGISTERS_3_13_port
                           , S => n704, Z => n4061);
   U4614 : MUX2_X1 port map( A => REGISTERS_0_13_port, B => REGISTERS_2_13_port
                           , S => n704, Z => n4062);
   U4615 : MUX2_X1 port map( A => n4062, B => n4061, S => n744, Z => n4063);
   U4616 : MUX2_X1 port map( A => n4063, B => n4060, S => n674, Z => n4064);
   U4617 : MUX2_X1 port map( A => n4064, B => n4057, S => r3007_A_3_port, Z => 
                           n4065);
   U4618 : MUX2_X1 port map( A => n4065, B => n4050, S => r3007_A_4_port, Z => 
                           n4066);
   U4619 : MUX2_X1 port map( A => n4066, B => n4035, S => ADD_RD1_5_port, Z => 
                           N4407);
   U4620 : MUX2_X1 port map( A => REGISTERS_37_14_port, B => 
                           REGISTERS_39_14_port, S => n704, Z => n4067);
   U4621 : MUX2_X1 port map( A => REGISTERS_36_14_port, B => 
                           REGISTERS_38_14_port, S => n704, Z => n4068);
   U4622 : MUX2_X1 port map( A => n4068, B => n4067, S => n744, Z => n4069);
   U4623 : MUX2_X1 port map( A => REGISTERS_33_14_port, B => 
                           REGISTERS_35_14_port, S => n703, Z => n4070);
   U4624 : MUX2_X1 port map( A => REGISTERS_32_14_port, B => 
                           REGISTERS_34_14_port, S => n703, Z => n4071);
   U4625 : MUX2_X1 port map( A => n4071, B => n4070, S => n744, Z => n4072);
   U4626 : MUX2_X1 port map( A => n4072, B => n4069, S => n674, Z => n4073);
   U4627 : MUX2_X1 port map( A => REGISTERS_29_14_port, B => 
                           REGISTERS_31_14_port, S => n703, Z => n4074);
   U4628 : MUX2_X1 port map( A => REGISTERS_28_14_port, B => 
                           REGISTERS_30_14_port, S => n703, Z => n4075);
   U4629 : MUX2_X1 port map( A => n4075, B => n4074, S => n743, Z => n4076);
   U4630 : MUX2_X1 port map( A => REGISTERS_25_14_port, B => 
                           REGISTERS_27_14_port, S => n703, Z => n4077);
   U4631 : MUX2_X1 port map( A => REGISTERS_24_14_port, B => 
                           REGISTERS_26_14_port, S => n703, Z => n4078);
   U4632 : MUX2_X1 port map( A => n4078, B => n4077, S => n743, Z => n4079);
   U4633 : MUX2_X1 port map( A => n4079, B => n4076, S => n674, Z => n4080);
   U4634 : MUX2_X1 port map( A => REGISTERS_21_14_port, B => 
                           REGISTERS_23_14_port, S => n703, Z => n4081);
   U4635 : MUX2_X1 port map( A => REGISTERS_20_14_port, B => 
                           REGISTERS_22_14_port, S => n703, Z => n4082);
   U4636 : MUX2_X1 port map( A => n4082, B => n4081, S => n743, Z => n4083);
   U4637 : MUX2_X1 port map( A => REGISTERS_17_14_port, B => 
                           REGISTERS_19_14_port, S => n703, Z => n4084);
   U4638 : MUX2_X1 port map( A => REGISTERS_16_14_port, B => 
                           REGISTERS_18_14_port, S => n703, Z => n4085);
   U4639 : MUX2_X1 port map( A => n4085, B => n4084, S => n743, Z => n4086);
   U4640 : MUX2_X1 port map( A => n4086, B => n4083, S => n674, Z => n4087);
   U4641 : MUX2_X1 port map( A => n4087, B => n4080, S => r3007_A_3_port, Z => 
                           n4088);
   U4642 : MUX2_X1 port map( A => REGISTERS_13_14_port, B => 
                           REGISTERS_15_14_port, S => n703, Z => n4089);
   U4643 : MUX2_X1 port map( A => REGISTERS_12_14_port, B => 
                           REGISTERS_14_14_port, S => n703, Z => n4090);
   U4644 : MUX2_X1 port map( A => n4090, B => n4089, S => n743, Z => n4091);
   U4645 : MUX2_X1 port map( A => REGISTERS_9_14_port, B => 
                           REGISTERS_11_14_port, S => n703, Z => n4092);
   U4646 : MUX2_X1 port map( A => REGISTERS_8_14_port, B => 
                           REGISTERS_10_14_port, S => n703, Z => n4093);
   U4647 : MUX2_X1 port map( A => n4093, B => n4092, S => n743, Z => n4094);
   U4648 : MUX2_X1 port map( A => n4094, B => n4091, S => n674, Z => n4095);
   U4649 : MUX2_X1 port map( A => REGISTERS_5_14_port, B => REGISTERS_7_14_port
                           , S => n703, Z => n4096);
   U4650 : MUX2_X1 port map( A => REGISTERS_4_14_port, B => REGISTERS_6_14_port
                           , S => n702, Z => n4097);
   U4651 : MUX2_X1 port map( A => n4097, B => n4096, S => n743, Z => n4098);
   U4652 : MUX2_X1 port map( A => REGISTERS_1_14_port, B => REGISTERS_3_14_port
                           , S => n702, Z => n4099);
   U4653 : MUX2_X1 port map( A => REGISTERS_0_14_port, B => REGISTERS_2_14_port
                           , S => n702, Z => n4100);
   U4654 : MUX2_X1 port map( A => n4100, B => n4099, S => n743, Z => n4101);
   U4655 : MUX2_X1 port map( A => n4101, B => n4098, S => n674, Z => n4102);
   U4656 : MUX2_X1 port map( A => n4102, B => n4095, S => r3007_A_3_port, Z => 
                           n4103);
   U4657 : MUX2_X1 port map( A => n4103, B => n4088, S => r3007_A_4_port, Z => 
                           n4104);
   U4658 : MUX2_X1 port map( A => n4104, B => n4073, S => ADD_RD1_5_port, Z => 
                           N4406);
   U4659 : MUX2_X1 port map( A => REGISTERS_37_15_port, B => 
                           REGISTERS_39_15_port, S => n702, Z => n4105);
   U4660 : MUX2_X1 port map( A => REGISTERS_36_15_port, B => 
                           REGISTERS_38_15_port, S => n702, Z => n4106);
   U4661 : MUX2_X1 port map( A => n4106, B => n4105, S => n743, Z => n4107);
   U4662 : MUX2_X1 port map( A => REGISTERS_33_15_port, B => 
                           REGISTERS_35_15_port, S => n702, Z => n4108);
   U4663 : MUX2_X1 port map( A => REGISTERS_32_15_port, B => 
                           REGISTERS_34_15_port, S => n702, Z => n4109);
   U4664 : MUX2_X1 port map( A => n4109, B => n4108, S => n743, Z => n4110);
   U4665 : MUX2_X1 port map( A => n4110, B => n4107, S => n674, Z => n4111);
   U4666 : MUX2_X1 port map( A => REGISTERS_29_15_port, B => 
                           REGISTERS_31_15_port, S => n702, Z => n4112);
   U4667 : MUX2_X1 port map( A => REGISTERS_28_15_port, B => 
                           REGISTERS_30_15_port, S => n702, Z => n4113);
   U4668 : MUX2_X1 port map( A => n4113, B => n4112, S => n743, Z => n4114);
   U4669 : MUX2_X1 port map( A => REGISTERS_25_15_port, B => 
                           REGISTERS_27_15_port, S => n702, Z => n4115);
   U4670 : MUX2_X1 port map( A => REGISTERS_24_15_port, B => 
                           REGISTERS_26_15_port, S => n702, Z => n4116);
   U4671 : MUX2_X1 port map( A => n4116, B => n4115, S => n743, Z => n4117);
   U4672 : MUX2_X1 port map( A => n4117, B => n4114, S => n674, Z => n4118);
   U4673 : MUX2_X1 port map( A => REGISTERS_21_15_port, B => 
                           REGISTERS_23_15_port, S => n702, Z => n4119);
   U4674 : MUX2_X1 port map( A => REGISTERS_20_15_port, B => 
                           REGISTERS_22_15_port, S => n702, Z => n4120);
   U4675 : MUX2_X1 port map( A => n4120, B => n4119, S => n743, Z => n4121);
   U4676 : MUX2_X1 port map( A => REGISTERS_17_15_port, B => 
                           REGISTERS_19_15_port, S => n702, Z => n4122);
   U4677 : MUX2_X1 port map( A => REGISTERS_16_15_port, B => 
                           REGISTERS_18_15_port, S => n702, Z => n4123);
   U4678 : MUX2_X1 port map( A => n4123, B => n4122, S => n743, Z => n4124);
   U4679 : MUX2_X1 port map( A => n4124, B => n4121, S => n673, Z => n4125);
   U4680 : MUX2_X1 port map( A => n4125, B => n4118, S => r3007_A_3_port, Z => 
                           n4126);
   U4681 : MUX2_X1 port map( A => REGISTERS_13_15_port, B => 
                           REGISTERS_15_15_port, S => n701, Z => n4127);
   U4682 : MUX2_X1 port map( A => REGISTERS_12_15_port, B => 
                           REGISTERS_14_15_port, S => n701, Z => n4128);
   U4683 : MUX2_X1 port map( A => n4128, B => n4127, S => n743, Z => n4129);
   U4684 : MUX2_X1 port map( A => REGISTERS_9_15_port, B => 
                           REGISTERS_11_15_port, S => n701, Z => n4130);
   U4685 : MUX2_X1 port map( A => REGISTERS_8_15_port, B => 
                           REGISTERS_10_15_port, S => n701, Z => n4131);
   U4686 : MUX2_X1 port map( A => n4131, B => n4130, S => n742, Z => n4132);
   U4687 : MUX2_X1 port map( A => n4132, B => n4129, S => n673, Z => n4133);
   U4688 : MUX2_X1 port map( A => REGISTERS_5_15_port, B => REGISTERS_7_15_port
                           , S => n701, Z => n4134);
   U4689 : MUX2_X1 port map( A => REGISTERS_4_15_port, B => REGISTERS_6_15_port
                           , S => n701, Z => n4135);
   U4690 : MUX2_X1 port map( A => n4135, B => n4134, S => n742, Z => n4136);
   U4691 : MUX2_X1 port map( A => REGISTERS_1_15_port, B => REGISTERS_3_15_port
                           , S => n701, Z => n4137);
   U4692 : MUX2_X1 port map( A => REGISTERS_0_15_port, B => REGISTERS_2_15_port
                           , S => n701, Z => n4138);
   U4693 : MUX2_X1 port map( A => n4138, B => n4137, S => n742, Z => n4139);
   U4694 : MUX2_X1 port map( A => n4139, B => n4136, S => n673, Z => n4140);
   U4695 : MUX2_X1 port map( A => n4140, B => n4133, S => r3007_A_3_port, Z => 
                           n4141);
   U4696 : MUX2_X1 port map( A => n4141, B => n4126, S => r3007_A_4_port, Z => 
                           n4142);
   U4697 : MUX2_X1 port map( A => n4142, B => n4111, S => ADD_RD1_5_port, Z => 
                           N4405);
   U4698 : MUX2_X1 port map( A => REGISTERS_37_16_port, B => 
                           REGISTERS_39_16_port, S => n701, Z => n4143);
   U4699 : MUX2_X1 port map( A => REGISTERS_36_16_port, B => 
                           REGISTERS_38_16_port, S => n701, Z => n4144);
   U4700 : MUX2_X1 port map( A => n4144, B => n4143, S => n742, Z => n4145);
   U4701 : MUX2_X1 port map( A => REGISTERS_33_16_port, B => 
                           REGISTERS_35_16_port, S => n701, Z => n4146);
   U4702 : MUX2_X1 port map( A => REGISTERS_32_16_port, B => 
                           REGISTERS_34_16_port, S => n701, Z => n4147);
   U4703 : MUX2_X1 port map( A => n4147, B => n4146, S => n742, Z => n4148);
   U4704 : MUX2_X1 port map( A => n4148, B => n4145, S => n673, Z => n4149);
   U4705 : MUX2_X1 port map( A => REGISTERS_29_16_port, B => 
                           REGISTERS_31_16_port, S => n701, Z => n4150);
   U4706 : MUX2_X1 port map( A => REGISTERS_28_16_port, B => 
                           REGISTERS_30_16_port, S => n701, Z => n4151);
   U4707 : MUX2_X1 port map( A => n4151, B => n4150, S => n742, Z => n4152);
   U4708 : MUX2_X1 port map( A => REGISTERS_25_16_port, B => 
                           REGISTERS_27_16_port, S => n701, Z => n4153);
   U4709 : MUX2_X1 port map( A => REGISTERS_24_16_port, B => 
                           REGISTERS_26_16_port, S => n700, Z => n4154);
   U4710 : MUX2_X1 port map( A => n4154, B => n4153, S => n742, Z => n4155);
   U4711 : MUX2_X1 port map( A => n4155, B => n4152, S => n673, Z => n4156);
   U4712 : MUX2_X1 port map( A => REGISTERS_21_16_port, B => 
                           REGISTERS_23_16_port, S => n700, Z => n4157);
   U4713 : MUX2_X1 port map( A => REGISTERS_20_16_port, B => 
                           REGISTERS_22_16_port, S => n700, Z => n4158);
   U4714 : MUX2_X1 port map( A => n4158, B => n4157, S => n742, Z => n4159);
   U4715 : MUX2_X1 port map( A => REGISTERS_17_16_port, B => 
                           REGISTERS_19_16_port, S => n700, Z => n4160);
   U4716 : MUX2_X1 port map( A => REGISTERS_16_16_port, B => 
                           REGISTERS_18_16_port, S => n700, Z => n4161);
   U4717 : MUX2_X1 port map( A => n4161, B => n4160, S => n742, Z => n4162);
   U4718 : MUX2_X1 port map( A => n4162, B => n4159, S => n673, Z => n4163);
   U4719 : MUX2_X1 port map( A => n4163, B => n4156, S => r3007_A_3_port, Z => 
                           n4164);
   U4720 : MUX2_X1 port map( A => REGISTERS_13_16_port, B => 
                           REGISTERS_15_16_port, S => n700, Z => n4165);
   U4721 : MUX2_X1 port map( A => REGISTERS_12_16_port, B => 
                           REGISTERS_14_16_port, S => n700, Z => n4166);
   U4722 : MUX2_X1 port map( A => n4166, B => n4165, S => n742, Z => n4167);
   U4723 : MUX2_X1 port map( A => REGISTERS_9_16_port, B => 
                           REGISTERS_11_16_port, S => n700, Z => n4168);
   U4724 : MUX2_X1 port map( A => REGISTERS_8_16_port, B => 
                           REGISTERS_10_16_port, S => n700, Z => n4169);
   U4725 : MUX2_X1 port map( A => n4169, B => n4168, S => n742, Z => n4170);
   U4726 : MUX2_X1 port map( A => n4170, B => n4167, S => n673, Z => n4171);
   U4727 : MUX2_X1 port map( A => REGISTERS_5_16_port, B => REGISTERS_7_16_port
                           , S => n700, Z => n4172);
   U4728 : MUX2_X1 port map( A => REGISTERS_4_16_port, B => REGISTERS_6_16_port
                           , S => n700, Z => n4173);
   U4729 : MUX2_X1 port map( A => n4173, B => n4172, S => n742, Z => n4174);
   U4730 : MUX2_X1 port map( A => REGISTERS_1_16_port, B => REGISTERS_3_16_port
                           , S => n700, Z => n4175);
   U4731 : MUX2_X1 port map( A => REGISTERS_0_16_port, B => REGISTERS_2_16_port
                           , S => n700, Z => n4176);
   U4732 : MUX2_X1 port map( A => n4176, B => n4175, S => n742, Z => n4177);
   U4733 : MUX2_X1 port map( A => n4177, B => n4174, S => n673, Z => n4178);
   U4734 : MUX2_X1 port map( A => n4178, B => n4171, S => r3007_A_3_port, Z => 
                           n4179);
   U4735 : MUX2_X1 port map( A => n4179, B => n4164, S => r3007_A_4_port, Z => 
                           n4180);
   U4736 : MUX2_X1 port map( A => n4180, B => n4149, S => ADD_RD1_5_port, Z => 
                           N4404);
   U4737 : MUX2_X1 port map( A => REGISTERS_37_17_port, B => 
                           REGISTERS_39_17_port, S => n700, Z => n4181);
   U4738 : MUX2_X1 port map( A => REGISTERS_36_17_port, B => 
                           REGISTERS_38_17_port, S => n700, Z => n4182);
   U4739 : MUX2_X1 port map( A => n4182, B => n4181, S => n742, Z => n4183);
   U4740 : MUX2_X1 port map( A => REGISTERS_33_17_port, B => 
                           REGISTERS_35_17_port, S => n699, Z => n4184);
   U4741 : MUX2_X1 port map( A => REGISTERS_32_17_port, B => 
                           REGISTERS_34_17_port, S => n699, Z => n4185);
   U4742 : MUX2_X1 port map( A => n4185, B => n4184, S => n742, Z => n4186);
   U4743 : MUX2_X1 port map( A => n4186, B => n4183, S => n673, Z => n4187);
   U4744 : MUX2_X1 port map( A => REGISTERS_29_17_port, B => 
                           REGISTERS_31_17_port, S => n699, Z => n4188);
   U4745 : MUX2_X1 port map( A => REGISTERS_28_17_port, B => 
                           REGISTERS_30_17_port, S => n699, Z => n4189);
   U4746 : MUX2_X1 port map( A => n4189, B => n4188, S => n741, Z => n4190);
   U4747 : MUX2_X1 port map( A => REGISTERS_25_17_port, B => 
                           REGISTERS_27_17_port, S => n699, Z => n4191);
   U4748 : MUX2_X1 port map( A => REGISTERS_24_17_port, B => 
                           REGISTERS_26_17_port, S => n699, Z => n4192);
   U4749 : MUX2_X1 port map( A => n4192, B => n4191, S => n741, Z => n4193);
   U4750 : MUX2_X1 port map( A => n4193, B => n4190, S => n673, Z => n4194);
   U4751 : MUX2_X1 port map( A => REGISTERS_21_17_port, B => 
                           REGISTERS_23_17_port, S => n699, Z => n4195);
   U4752 : MUX2_X1 port map( A => REGISTERS_20_17_port, B => 
                           REGISTERS_22_17_port, S => n699, Z => n4196);
   U4753 : MUX2_X1 port map( A => n4196, B => n4195, S => n741, Z => n4197);
   U4754 : MUX2_X1 port map( A => REGISTERS_17_17_port, B => 
                           REGISTERS_19_17_port, S => n699, Z => n4198);
   U4755 : MUX2_X1 port map( A => REGISTERS_16_17_port, B => 
                           REGISTERS_18_17_port, S => n699, Z => n4199);
   U4756 : MUX2_X1 port map( A => n4199, B => n4198, S => n741, Z => n4200);
   U4757 : MUX2_X1 port map( A => n4200, B => n4197, S => n673, Z => n4201);
   U4758 : MUX2_X1 port map( A => n4201, B => n4194, S => r3007_A_3_port, Z => 
                           n4202);
   U4759 : MUX2_X1 port map( A => REGISTERS_13_17_port, B => 
                           REGISTERS_15_17_port, S => n699, Z => n4203);
   U4760 : MUX2_X1 port map( A => REGISTERS_12_17_port, B => 
                           REGISTERS_14_17_port, S => n699, Z => n4204);
   U4761 : MUX2_X1 port map( A => n4204, B => n4203, S => n741, Z => n4205);
   U4762 : MUX2_X1 port map( A => REGISTERS_9_17_port, B => 
                           REGISTERS_11_17_port, S => n699, Z => n4206);
   U4763 : MUX2_X1 port map( A => REGISTERS_8_17_port, B => 
                           REGISTERS_10_17_port, S => n699, Z => n4207);
   U4764 : MUX2_X1 port map( A => n4207, B => n4206, S => n741, Z => n4208);
   U4765 : MUX2_X1 port map( A => n4208, B => n4205, S => n673, Z => n4209);
   U4766 : MUX2_X1 port map( A => REGISTERS_5_17_port, B => REGISTERS_7_17_port
                           , S => n699, Z => n4210);
   U4767 : MUX2_X1 port map( A => REGISTERS_4_17_port, B => REGISTERS_6_17_port
                           , S => n698, Z => n4211);
   U4768 : MUX2_X1 port map( A => n4211, B => n4210, S => n741, Z => n4212);
   U4769 : MUX2_X1 port map( A => REGISTERS_1_17_port, B => REGISTERS_3_17_port
                           , S => n698, Z => n4213);
   U4770 : MUX2_X1 port map( A => REGISTERS_0_17_port, B => REGISTERS_2_17_port
                           , S => n698, Z => n4214);
   U4771 : MUX2_X1 port map( A => n4214, B => n4213, S => n741, Z => n4215);
   U4772 : MUX2_X1 port map( A => n4215, B => n4212, S => n673, Z => n4216);
   U4773 : MUX2_X1 port map( A => n4216, B => n4209, S => r3007_A_3_port, Z => 
                           n4217);
   U4774 : MUX2_X1 port map( A => n4217, B => n4202, S => r3007_A_4_port, Z => 
                           n4218);
   U4775 : MUX2_X1 port map( A => n4218, B => n4187, S => ADD_RD1_5_port, Z => 
                           N4403);
   U4776 : MUX2_X1 port map( A => REGISTERS_37_18_port, B => 
                           REGISTERS_39_18_port, S => n698, Z => n4219);
   U4777 : MUX2_X1 port map( A => REGISTERS_36_18_port, B => 
                           REGISTERS_38_18_port, S => n698, Z => n4220);
   U4778 : MUX2_X1 port map( A => n4220, B => n4219, S => n741, Z => n4221);
   U4779 : MUX2_X1 port map( A => REGISTERS_33_18_port, B => 
                           REGISTERS_35_18_port, S => n698, Z => n4222);
   U4780 : MUX2_X1 port map( A => REGISTERS_32_18_port, B => 
                           REGISTERS_34_18_port, S => n698, Z => n4223);
   U4781 : MUX2_X1 port map( A => n4223, B => n4222, S => n741, Z => n4224);
   U4782 : MUX2_X1 port map( A => n4224, B => n4221, S => n673, Z => n4225);
   U4783 : MUX2_X1 port map( A => REGISTERS_29_18_port, B => 
                           REGISTERS_31_18_port, S => n698, Z => n4226);
   U4784 : MUX2_X1 port map( A => REGISTERS_28_18_port, B => 
                           REGISTERS_30_18_port, S => n698, Z => n4227);
   U4785 : MUX2_X1 port map( A => n4227, B => n4226, S => n741, Z => n4228);
   U4786 : MUX2_X1 port map( A => REGISTERS_25_18_port, B => 
                           REGISTERS_27_18_port, S => n698, Z => n4229);
   U4787 : MUX2_X1 port map( A => REGISTERS_24_18_port, B => 
                           REGISTERS_26_18_port, S => n698, Z => n4230);
   U4788 : MUX2_X1 port map( A => n4230, B => n4229, S => n741, Z => n4231);
   U4789 : MUX2_X1 port map( A => n4231, B => n4228, S => n672, Z => n4232);
   U4790 : MUX2_X1 port map( A => REGISTERS_21_18_port, B => 
                           REGISTERS_23_18_port, S => n698, Z => n4233);
   U4791 : MUX2_X1 port map( A => REGISTERS_20_18_port, B => 
                           REGISTERS_22_18_port, S => n698, Z => n4234);
   U4792 : MUX2_X1 port map( A => n4234, B => n4233, S => n741, Z => n4235);
   U4793 : MUX2_X1 port map( A => REGISTERS_17_18_port, B => 
                           REGISTERS_19_18_port, S => n698, Z => n4236);
   U4794 : MUX2_X1 port map( A => REGISTERS_16_18_port, B => 
                           REGISTERS_18_18_port, S => n698, Z => n4237);
   U4795 : MUX2_X1 port map( A => n4237, B => n4236, S => n741, Z => n4238);
   U4796 : MUX2_X1 port map( A => n4238, B => n4235, S => n672, Z => n4239);
   U4797 : MUX2_X1 port map( A => n4239, B => n4232, S => r3007_A_3_port, Z => 
                           n4240);
   U4798 : MUX2_X1 port map( A => REGISTERS_13_18_port, B => 
                           REGISTERS_15_18_port, S => n697, Z => n4241);
   U4799 : MUX2_X1 port map( A => REGISTERS_12_18_port, B => 
                           REGISTERS_14_18_port, S => n697, Z => n4242);
   U4800 : MUX2_X1 port map( A => n4242, B => n4241, S => n741, Z => n4243);
   U4801 : MUX2_X1 port map( A => REGISTERS_9_18_port, B => 
                           REGISTERS_11_18_port, S => n697, Z => n4244);
   U4802 : MUX2_X1 port map( A => REGISTERS_8_18_port, B => 
                           REGISTERS_10_18_port, S => n697, Z => n4245);
   U4803 : MUX2_X1 port map( A => n4245, B => n4244, S => n740, Z => n4246);
   U4804 : MUX2_X1 port map( A => n4246, B => n4243, S => n672, Z => n4247);
   U4805 : MUX2_X1 port map( A => REGISTERS_5_18_port, B => REGISTERS_7_18_port
                           , S => n697, Z => n4248);
   U4806 : MUX2_X1 port map( A => REGISTERS_4_18_port, B => REGISTERS_6_18_port
                           , S => n697, Z => n4249);
   U4807 : MUX2_X1 port map( A => n4249, B => n4248, S => n740, Z => n4250);
   U4808 : MUX2_X1 port map( A => REGISTERS_1_18_port, B => REGISTERS_3_18_port
                           , S => n697, Z => n4251);
   U4809 : MUX2_X1 port map( A => REGISTERS_0_18_port, B => REGISTERS_2_18_port
                           , S => n697, Z => n4252);
   U4810 : MUX2_X1 port map( A => n4252, B => n4251, S => n740, Z => n4253);
   U4811 : MUX2_X1 port map( A => n4253, B => n4250, S => n672, Z => n4254);
   U4812 : MUX2_X1 port map( A => n4254, B => n4247, S => r3007_A_3_port, Z => 
                           n4255);
   U4813 : MUX2_X1 port map( A => n4255, B => n4240, S => r3007_A_4_port, Z => 
                           n4256);
   U4814 : MUX2_X1 port map( A => n4256, B => n4225, S => ADD_RD1_5_port, Z => 
                           N4402);
   U4815 : MUX2_X1 port map( A => REGISTERS_37_19_port, B => 
                           REGISTERS_39_19_port, S => n697, Z => n4257);
   U4816 : MUX2_X1 port map( A => REGISTERS_36_19_port, B => 
                           REGISTERS_38_19_port, S => n697, Z => n4258);
   U4817 : MUX2_X1 port map( A => n4258, B => n4257, S => n740, Z => n4259);
   U4818 : MUX2_X1 port map( A => REGISTERS_33_19_port, B => 
                           REGISTERS_35_19_port, S => n697, Z => n4260);
   U4819 : MUX2_X1 port map( A => REGISTERS_32_19_port, B => 
                           REGISTERS_34_19_port, S => n697, Z => n4261);
   U4820 : MUX2_X1 port map( A => n4261, B => n4260, S => n740, Z => n4262);
   U4821 : MUX2_X1 port map( A => n4262, B => n4259, S => n672, Z => n4263);
   U4822 : MUX2_X1 port map( A => REGISTERS_29_19_port, B => 
                           REGISTERS_31_19_port, S => n697, Z => n4264);
   U4823 : MUX2_X1 port map( A => REGISTERS_28_19_port, B => 
                           REGISTERS_30_19_port, S => n697, Z => n4265);
   U4824 : MUX2_X1 port map( A => n4265, B => n4264, S => n740, Z => n4266);
   U4825 : MUX2_X1 port map( A => REGISTERS_25_19_port, B => 
                           REGISTERS_27_19_port, S => n697, Z => n4267);
   U4826 : MUX2_X1 port map( A => REGISTERS_24_19_port, B => 
                           REGISTERS_26_19_port, S => n696, Z => n4268);
   U4827 : MUX2_X1 port map( A => n4268, B => n4267, S => n740, Z => n4269);
   U4828 : MUX2_X1 port map( A => n4269, B => n4266, S => n672, Z => n4270);
   U4829 : MUX2_X1 port map( A => REGISTERS_21_19_port, B => 
                           REGISTERS_23_19_port, S => n696, Z => n4271);
   U4830 : MUX2_X1 port map( A => REGISTERS_20_19_port, B => 
                           REGISTERS_22_19_port, S => n696, Z => n4272);
   U4831 : MUX2_X1 port map( A => n4272, B => n4271, S => n740, Z => n4273);
   U4832 : MUX2_X1 port map( A => REGISTERS_17_19_port, B => 
                           REGISTERS_19_19_port, S => n696, Z => n4274);
   U4833 : MUX2_X1 port map( A => REGISTERS_16_19_port, B => 
                           REGISTERS_18_19_port, S => n696, Z => n4275);
   U4834 : MUX2_X1 port map( A => n4275, B => n4274, S => n740, Z => n4276);
   U4835 : MUX2_X1 port map( A => n4276, B => n4273, S => n672, Z => n4277);
   U4836 : MUX2_X1 port map( A => n4277, B => n4270, S => r3007_A_3_port, Z => 
                           n4278);
   U4837 : MUX2_X1 port map( A => REGISTERS_13_19_port, B => 
                           REGISTERS_15_19_port, S => n696, Z => n4279);
   U4838 : MUX2_X1 port map( A => REGISTERS_12_19_port, B => 
                           REGISTERS_14_19_port, S => n696, Z => n4280);
   U4839 : MUX2_X1 port map( A => n4280, B => n4279, S => n740, Z => n4281);
   U4840 : MUX2_X1 port map( A => REGISTERS_9_19_port, B => 
                           REGISTERS_11_19_port, S => n696, Z => n4282);
   U4841 : MUX2_X1 port map( A => REGISTERS_8_19_port, B => 
                           REGISTERS_10_19_port, S => n696, Z => n4283);
   U4842 : MUX2_X1 port map( A => n4283, B => n4282, S => n740, Z => n4284);
   U4843 : MUX2_X1 port map( A => n4284, B => n4281, S => n672, Z => n4285);
   U4844 : MUX2_X1 port map( A => REGISTERS_5_19_port, B => REGISTERS_7_19_port
                           , S => n696, Z => n4286);
   U4845 : MUX2_X1 port map( A => REGISTERS_4_19_port, B => REGISTERS_6_19_port
                           , S => n696, Z => n4287);
   U4846 : MUX2_X1 port map( A => n4287, B => n4286, S => n740, Z => n4288);
   U4847 : MUX2_X1 port map( A => REGISTERS_1_19_port, B => REGISTERS_3_19_port
                           , S => n696, Z => n4289);
   U4848 : MUX2_X1 port map( A => REGISTERS_0_19_port, B => REGISTERS_2_19_port
                           , S => n696, Z => n4290);
   U4849 : MUX2_X1 port map( A => n4290, B => n4289, S => n740, Z => n4291);
   U4850 : MUX2_X1 port map( A => n4291, B => n4288, S => n672, Z => n4292);
   U4851 : MUX2_X1 port map( A => n4292, B => n4285, S => r3007_A_3_port, Z => 
                           n4293);
   U4852 : MUX2_X1 port map( A => n4293, B => n4278, S => r3007_A_4_port, Z => 
                           n4294);
   U4853 : MUX2_X1 port map( A => n4294, B => n4263, S => ADD_RD1_5_port, Z => 
                           N4401);
   U4854 : MUX2_X1 port map( A => REGISTERS_37_20_port, B => 
                           REGISTERS_39_20_port, S => n696, Z => n4295);
   U4855 : MUX2_X1 port map( A => REGISTERS_36_20_port, B => 
                           REGISTERS_38_20_port, S => n696, Z => n4296);
   U4856 : MUX2_X1 port map( A => n4296, B => n4295, S => n740, Z => n4297);
   U4857 : MUX2_X1 port map( A => REGISTERS_33_20_port, B => 
                           REGISTERS_35_20_port, S => n695, Z => n4298);
   U4858 : MUX2_X1 port map( A => REGISTERS_32_20_port, B => 
                           REGISTERS_34_20_port, S => n695, Z => n4299);
   U4859 : MUX2_X1 port map( A => n4299, B => n4298, S => n740, Z => n4300);
   U4860 : MUX2_X1 port map( A => n4300, B => n4297, S => n672, Z => n4301);
   U4861 : MUX2_X1 port map( A => REGISTERS_29_20_port, B => 
                           REGISTERS_31_20_port, S => n695, Z => n4302);
   U4862 : MUX2_X1 port map( A => REGISTERS_28_20_port, B => 
                           REGISTERS_30_20_port, S => n695, Z => n4303);
   U4863 : MUX2_X1 port map( A => n4303, B => n4302, S => n739, Z => n4304);
   U4864 : MUX2_X1 port map( A => REGISTERS_25_20_port, B => 
                           REGISTERS_27_20_port, S => n695, Z => n4305);
   U4865 : MUX2_X1 port map( A => REGISTERS_24_20_port, B => 
                           REGISTERS_26_20_port, S => n695, Z => n4306);
   U4866 : MUX2_X1 port map( A => n4306, B => n4305, S => n739, Z => n4307);
   U4867 : MUX2_X1 port map( A => n4307, B => n4304, S => n672, Z => n4308);
   U4868 : MUX2_X1 port map( A => REGISTERS_21_20_port, B => 
                           REGISTERS_23_20_port, S => n695, Z => n4309);
   U4869 : MUX2_X1 port map( A => REGISTERS_20_20_port, B => 
                           REGISTERS_22_20_port, S => n695, Z => n4310);
   U4870 : MUX2_X1 port map( A => n4310, B => n4309, S => n739, Z => n4311);
   U4871 : MUX2_X1 port map( A => REGISTERS_17_20_port, B => 
                           REGISTERS_19_20_port, S => n695, Z => n4312);
   U4872 : MUX2_X1 port map( A => REGISTERS_16_20_port, B => 
                           REGISTERS_18_20_port, S => n695, Z => n4313);
   U4873 : MUX2_X1 port map( A => n4313, B => n4312, S => n739, Z => n4314);
   U4874 : MUX2_X1 port map( A => n4314, B => n4311, S => n672, Z => n4315);
   U4875 : MUX2_X1 port map( A => n4315, B => n4308, S => r3007_A_3_port, Z => 
                           n4316);
   U4876 : MUX2_X1 port map( A => REGISTERS_13_20_port, B => 
                           REGISTERS_15_20_port, S => n695, Z => n4317);
   U4877 : MUX2_X1 port map( A => REGISTERS_12_20_port, B => 
                           REGISTERS_14_20_port, S => n695, Z => n4318);
   U4878 : MUX2_X1 port map( A => n4318, B => n4317, S => n739, Z => n4319);
   U4879 : MUX2_X1 port map( A => REGISTERS_9_20_port, B => 
                           REGISTERS_11_20_port, S => n695, Z => n4320);
   U4880 : MUX2_X1 port map( A => REGISTERS_8_20_port, B => 
                           REGISTERS_10_20_port, S => n695, Z => n4321);
   U4881 : MUX2_X1 port map( A => n4321, B => n4320, S => n739, Z => n4322);
   U4882 : MUX2_X1 port map( A => n4322, B => n4319, S => n672, Z => n4323);
   U4883 : MUX2_X1 port map( A => REGISTERS_5_20_port, B => REGISTERS_7_20_port
                           , S => n695, Z => n4324);
   U4884 : MUX2_X1 port map( A => REGISTERS_4_20_port, B => REGISTERS_6_20_port
                           , S => n694, Z => n4325);
   U4885 : MUX2_X1 port map( A => n4325, B => n4324, S => n739, Z => n4326);
   U4886 : MUX2_X1 port map( A => REGISTERS_1_20_port, B => REGISTERS_3_20_port
                           , S => n694, Z => n4327);
   U4887 : MUX2_X1 port map( A => REGISTERS_0_20_port, B => REGISTERS_2_20_port
                           , S => n694, Z => n4328);
   U4888 : MUX2_X1 port map( A => n4328, B => n4327, S => n739, Z => n4329);
   U4889 : MUX2_X1 port map( A => n4329, B => n4326, S => n672, Z => n4330);
   U4890 : MUX2_X1 port map( A => n4330, B => n4323, S => r3007_A_3_port, Z => 
                           n4331);
   U4891 : MUX2_X1 port map( A => n4331, B => n4316, S => r3007_A_4_port, Z => 
                           n4332);
   U4892 : MUX2_X1 port map( A => n4332, B => n4301, S => ADD_RD1_5_port, Z => 
                           N4400);
   U4893 : MUX2_X1 port map( A => REGISTERS_37_21_port, B => 
                           REGISTERS_39_21_port, S => n694, Z => n4333);
   U4894 : MUX2_X1 port map( A => REGISTERS_36_21_port, B => 
                           REGISTERS_38_21_port, S => n694, Z => n4334);
   U4895 : MUX2_X1 port map( A => n4334, B => n4333, S => n739, Z => n4335);
   U4896 : MUX2_X1 port map( A => REGISTERS_33_21_port, B => 
                           REGISTERS_35_21_port, S => n694, Z => n4336);
   U4897 : MUX2_X1 port map( A => REGISTERS_32_21_port, B => 
                           REGISTERS_34_21_port, S => n694, Z => n4337);
   U4898 : MUX2_X1 port map( A => n4337, B => n4336, S => n739, Z => n4338);
   U4899 : MUX2_X1 port map( A => n4338, B => n4335, S => n671, Z => n4339);
   U4900 : MUX2_X1 port map( A => REGISTERS_29_21_port, B => 
                           REGISTERS_31_21_port, S => n694, Z => n4340);
   U4901 : MUX2_X1 port map( A => REGISTERS_28_21_port, B => 
                           REGISTERS_30_21_port, S => n694, Z => n4341);
   U4902 : MUX2_X1 port map( A => n4341, B => n4340, S => n739, Z => n4342);
   U4903 : MUX2_X1 port map( A => REGISTERS_25_21_port, B => 
                           REGISTERS_27_21_port, S => n694, Z => n4343);
   U4904 : MUX2_X1 port map( A => REGISTERS_24_21_port, B => 
                           REGISTERS_26_21_port, S => n694, Z => n4344);
   U4905 : MUX2_X1 port map( A => n4344, B => n4343, S => n739, Z => n4345);
   U4906 : MUX2_X1 port map( A => n4345, B => n4342, S => n671, Z => n4346);
   U4907 : MUX2_X1 port map( A => REGISTERS_21_21_port, B => 
                           REGISTERS_23_21_port, S => n694, Z => n4347);
   U4908 : MUX2_X1 port map( A => REGISTERS_20_21_port, B => 
                           REGISTERS_22_21_port, S => n694, Z => n4348);
   U4909 : MUX2_X1 port map( A => n4348, B => n4347, S => n739, Z => n4349);
   U4910 : MUX2_X1 port map( A => REGISTERS_17_21_port, B => 
                           REGISTERS_19_21_port, S => n694, Z => n4350);
   U4911 : MUX2_X1 port map( A => REGISTERS_16_21_port, B => 
                           REGISTERS_18_21_port, S => n694, Z => n4351);
   U4912 : MUX2_X1 port map( A => n4351, B => n4350, S => n739, Z => n4352);
   U4913 : MUX2_X1 port map( A => n4352, B => n4349, S => n671, Z => n4353);
   U4914 : MUX2_X1 port map( A => n4353, B => n4346, S => r3007_A_3_port, Z => 
                           n4354);
   U4915 : MUX2_X1 port map( A => REGISTERS_13_21_port, B => 
                           REGISTERS_15_21_port, S => n693, Z => n4355);
   U4916 : MUX2_X1 port map( A => REGISTERS_12_21_port, B => 
                           REGISTERS_14_21_port, S => n693, Z => n4356);
   U4917 : MUX2_X1 port map( A => n4356, B => n4355, S => n739, Z => n4357);
   U4918 : MUX2_X1 port map( A => REGISTERS_9_21_port, B => 
                           REGISTERS_11_21_port, S => n693, Z => n4358);
   U4919 : MUX2_X1 port map( A => REGISTERS_8_21_port, B => 
                           REGISTERS_10_21_port, S => n693, Z => n4359);
   U4920 : MUX2_X1 port map( A => n4359, B => n4358, S => n738, Z => n4360);
   U4921 : MUX2_X1 port map( A => n4360, B => n4357, S => n671, Z => n4361);
   U4922 : MUX2_X1 port map( A => REGISTERS_5_21_port, B => REGISTERS_7_21_port
                           , S => n693, Z => n4362);
   U4923 : MUX2_X1 port map( A => REGISTERS_4_21_port, B => REGISTERS_6_21_port
                           , S => n693, Z => n4363);
   U4924 : MUX2_X1 port map( A => n4363, B => n4362, S => n738, Z => n4364);
   U4925 : MUX2_X1 port map( A => REGISTERS_1_21_port, B => REGISTERS_3_21_port
                           , S => n693, Z => n4365);
   U4926 : MUX2_X1 port map( A => REGISTERS_0_21_port, B => REGISTERS_2_21_port
                           , S => n693, Z => n4366);
   U4927 : MUX2_X1 port map( A => n4366, B => n4365, S => n738, Z => n4367);
   U4928 : MUX2_X1 port map( A => n4367, B => n4364, S => n671, Z => n4368);
   U4929 : MUX2_X1 port map( A => n4368, B => n4361, S => r3007_A_3_port, Z => 
                           n4369);
   U4930 : MUX2_X1 port map( A => n4369, B => n4354, S => r3007_A_4_port, Z => 
                           n4370);
   U4931 : MUX2_X1 port map( A => n4370, B => n4339, S => ADD_RD1_5_port, Z => 
                           N4399);
   U4932 : MUX2_X1 port map( A => REGISTERS_37_22_port, B => 
                           REGISTERS_39_22_port, S => n693, Z => n4371);
   U4933 : MUX2_X1 port map( A => REGISTERS_36_22_port, B => 
                           REGISTERS_38_22_port, S => n693, Z => n4372);
   U4934 : MUX2_X1 port map( A => n4372, B => n4371, S => n738, Z => n4373);
   U4935 : MUX2_X1 port map( A => REGISTERS_33_22_port, B => 
                           REGISTERS_35_22_port, S => n693, Z => n4374);
   U4936 : MUX2_X1 port map( A => REGISTERS_32_22_port, B => 
                           REGISTERS_34_22_port, S => n693, Z => n4375);
   U4937 : MUX2_X1 port map( A => n4375, B => n4374, S => n738, Z => n4376);
   U4938 : MUX2_X1 port map( A => n4376, B => n4373, S => n671, Z => n4377);
   U4939 : MUX2_X1 port map( A => REGISTERS_29_22_port, B => 
                           REGISTERS_31_22_port, S => n693, Z => n4378);
   U4940 : MUX2_X1 port map( A => REGISTERS_28_22_port, B => 
                           REGISTERS_30_22_port, S => n693, Z => n4379);
   U4941 : MUX2_X1 port map( A => n4379, B => n4378, S => n738, Z => n4380);
   U4942 : MUX2_X1 port map( A => REGISTERS_25_22_port, B => 
                           REGISTERS_27_22_port, S => n693, Z => n4381);
   U4943 : MUX2_X1 port map( A => REGISTERS_24_22_port, B => 
                           REGISTERS_26_22_port, S => n692, Z => n4382);
   U4944 : MUX2_X1 port map( A => n4382, B => n4381, S => n738, Z => n4383);
   U4945 : MUX2_X1 port map( A => n4383, B => n4380, S => n671, Z => n4384);
   U4946 : MUX2_X1 port map( A => REGISTERS_21_22_port, B => 
                           REGISTERS_23_22_port, S => n692, Z => n4385);
   U4947 : MUX2_X1 port map( A => REGISTERS_20_22_port, B => 
                           REGISTERS_22_22_port, S => n692, Z => n4386);
   U4948 : MUX2_X1 port map( A => n4386, B => n4385, S => n738, Z => n4387);
   U4949 : MUX2_X1 port map( A => REGISTERS_17_22_port, B => 
                           REGISTERS_19_22_port, S => n692, Z => n4388);
   U4950 : MUX2_X1 port map( A => REGISTERS_16_22_port, B => 
                           REGISTERS_18_22_port, S => n692, Z => n4389_port);
   U4951 : MUX2_X1 port map( A => n4389_port, B => n4388, S => n738, Z => 
                           n4390_port);
   U4952 : MUX2_X1 port map( A => n4390_port, B => n4387, S => n671, Z => 
                           n4391_port);
   U4953 : MUX2_X1 port map( A => n4391_port, B => n4384, S => r3007_A_3_port, 
                           Z => n4392_port);
   U4954 : MUX2_X1 port map( A => REGISTERS_13_22_port, B => 
                           REGISTERS_15_22_port, S => n692, Z => n4393_port);
   U4955 : MUX2_X1 port map( A => REGISTERS_12_22_port, B => 
                           REGISTERS_14_22_port, S => n692, Z => n4394_port);
   U4956 : MUX2_X1 port map( A => n4394_port, B => n4393_port, S => n738, Z => 
                           n4395_port);
   U4957 : MUX2_X1 port map( A => REGISTERS_9_22_port, B => 
                           REGISTERS_11_22_port, S => n692, Z => n4396_port);
   U4958 : MUX2_X1 port map( A => REGISTERS_8_22_port, B => 
                           REGISTERS_10_22_port, S => n692, Z => n4397_port);
   U4959 : MUX2_X1 port map( A => n4397_port, B => n4396_port, S => n738, Z => 
                           n4398_port);
   U4960 : MUX2_X1 port map( A => n4398_port, B => n4395_port, S => n671, Z => 
                           n4399_port);
   U4961 : MUX2_X1 port map( A => REGISTERS_5_22_port, B => REGISTERS_7_22_port
                           , S => n692, Z => n4400_port);
   U4962 : MUX2_X1 port map( A => REGISTERS_4_22_port, B => REGISTERS_6_22_port
                           , S => n692, Z => n4401_port);
   U4963 : MUX2_X1 port map( A => n4401_port, B => n4400_port, S => n738, Z => 
                           n4402_port);
   U4964 : MUX2_X1 port map( A => REGISTERS_1_22_port, B => REGISTERS_3_22_port
                           , S => n692, Z => n4403_port);
   U4965 : MUX2_X1 port map( A => REGISTERS_0_22_port, B => REGISTERS_2_22_port
                           , S => n692, Z => n4404_port);
   U4966 : MUX2_X1 port map( A => n4404_port, B => n4403_port, S => n738, Z => 
                           n4405_port);
   U4967 : MUX2_X1 port map( A => n4405_port, B => n4402_port, S => n671, Z => 
                           n4406_port);
   U4968 : MUX2_X1 port map( A => n4406_port, B => n4399_port, S => 
                           r3007_A_3_port, Z => n4407_port);
   U4969 : MUX2_X1 port map( A => n4407_port, B => n4392_port, S => 
                           r3007_A_4_port, Z => n4408_port);
   U4970 : MUX2_X1 port map( A => n4408_port, B => n4377, S => ADD_RD1_5_port, 
                           Z => N4398);
   U4971 : MUX2_X1 port map( A => REGISTERS_37_23_port, B => 
                           REGISTERS_39_23_port, S => n692, Z => n4409_port);
   U4972 : MUX2_X1 port map( A => REGISTERS_36_23_port, B => 
                           REGISTERS_38_23_port, S => n692, Z => n4410_port);
   U4973 : MUX2_X1 port map( A => n4410_port, B => n4409_port, S => n738, Z => 
                           n4411_port);
   U4974 : MUX2_X1 port map( A => REGISTERS_33_23_port, B => 
                           REGISTERS_35_23_port, S => n691, Z => n4412_port);
   U4975 : MUX2_X1 port map( A => REGISTERS_32_23_port, B => 
                           REGISTERS_34_23_port, S => n691, Z => n4413_port);
   U4976 : MUX2_X1 port map( A => n4413_port, B => n4412_port, S => n738, Z => 
                           n4414_port);
   U4977 : MUX2_X1 port map( A => n4414_port, B => n4411_port, S => n671, Z => 
                           n4415_port);
   U4978 : MUX2_X1 port map( A => REGISTERS_29_23_port, B => 
                           REGISTERS_31_23_port, S => n691, Z => n4416_port);
   U4979 : MUX2_X1 port map( A => REGISTERS_28_23_port, B => 
                           REGISTERS_30_23_port, S => n691, Z => n4417_port);
   U4980 : MUX2_X1 port map( A => n4417_port, B => n4416_port, S => n737, Z => 
                           n4418_port);
   U4981 : MUX2_X1 port map( A => REGISTERS_25_23_port, B => 
                           REGISTERS_27_23_port, S => n691, Z => n4419_port);
   U4982 : MUX2_X1 port map( A => REGISTERS_24_23_port, B => 
                           REGISTERS_26_23_port, S => n691, Z => n4420_port);
   U4983 : MUX2_X1 port map( A => n4420_port, B => n4419_port, S => n737, Z => 
                           n4421);
   U4984 : MUX2_X1 port map( A => n4421, B => n4418_port, S => n671, Z => n4422
                           );
   U4985 : MUX2_X1 port map( A => REGISTERS_21_23_port, B => 
                           REGISTERS_23_23_port, S => n691, Z => n4423);
   U4986 : MUX2_X1 port map( A => REGISTERS_20_23_port, B => 
                           REGISTERS_22_23_port, S => n691, Z => n4424);
   U4987 : MUX2_X1 port map( A => n4424, B => n4423, S => n737, Z => n4425);
   U4988 : MUX2_X1 port map( A => REGISTERS_17_23_port, B => 
                           REGISTERS_19_23_port, S => n691, Z => n4426);
   U4989 : MUX2_X1 port map( A => REGISTERS_16_23_port, B => 
                           REGISTERS_18_23_port, S => n691, Z => n4427);
   U4990 : MUX2_X1 port map( A => n4427, B => n4426, S => n737, Z => n4428);
   U4991 : MUX2_X1 port map( A => n4428, B => n4425, S => n671, Z => n4429);
   U4992 : MUX2_X1 port map( A => n4429, B => n4422, S => r3007_A_3_port, Z => 
                           n4430);
   U4993 : MUX2_X1 port map( A => REGISTERS_13_23_port, B => 
                           REGISTERS_15_23_port, S => n691, Z => n4431);
   U4994 : MUX2_X1 port map( A => REGISTERS_12_23_port, B => 
                           REGISTERS_14_23_port, S => n691, Z => n4432);
   U4995 : MUX2_X1 port map( A => n4432, B => n4431, S => n737, Z => n4433);
   U4996 : MUX2_X1 port map( A => REGISTERS_9_23_port, B => 
                           REGISTERS_11_23_port, S => n691, Z => n4434);
   U4997 : MUX2_X1 port map( A => REGISTERS_8_23_port, B => 
                           REGISTERS_10_23_port, S => n691, Z => n4435);
   U4998 : MUX2_X1 port map( A => n4435, B => n4434, S => n737, Z => n4436);
   U4999 : MUX2_X1 port map( A => n4436, B => n4433, S => n671, Z => n4437);
   U5000 : MUX2_X1 port map( A => REGISTERS_5_23_port, B => REGISTERS_7_23_port
                           , S => n691, Z => n4438);
   U5001 : MUX2_X1 port map( A => REGISTERS_4_23_port, B => REGISTERS_6_23_port
                           , S => n690, Z => n4439);
   U5002 : MUX2_X1 port map( A => n4439, B => n4438, S => n737, Z => n4440);
   U5003 : MUX2_X1 port map( A => REGISTERS_1_23_port, B => REGISTERS_3_23_port
                           , S => n690, Z => n4441);
   U5004 : MUX2_X1 port map( A => REGISTERS_0_23_port, B => REGISTERS_2_23_port
                           , S => n690, Z => n4442);
   U5005 : MUX2_X1 port map( A => n4442, B => n4441, S => n737, Z => n4443);
   U5006 : MUX2_X1 port map( A => n4443, B => n4440, S => n670, Z => n4444);
   U5007 : MUX2_X1 port map( A => n4444, B => n4437, S => r3007_A_3_port, Z => 
                           n4445);
   U5008 : MUX2_X1 port map( A => n4445, B => n4430, S => r3007_A_4_port, Z => 
                           n4446);
   U5009 : MUX2_X1 port map( A => n4446, B => n4415_port, S => ADD_RD1_5_port, 
                           Z => N4397);
   U5010 : MUX2_X1 port map( A => REGISTERS_37_24_port, B => 
                           REGISTERS_39_24_port, S => n690, Z => n4447);
   U5011 : MUX2_X1 port map( A => REGISTERS_36_24_port, B => 
                           REGISTERS_38_24_port, S => n690, Z => n4448);
   U5012 : MUX2_X1 port map( A => n4448, B => n4447, S => n737, Z => n4449);
   U5013 : MUX2_X1 port map( A => REGISTERS_33_24_port, B => 
                           REGISTERS_35_24_port, S => n690, Z => n4450);
   U5014 : MUX2_X1 port map( A => REGISTERS_32_24_port, B => 
                           REGISTERS_34_24_port, S => n690, Z => n4451);
   U5015 : MUX2_X1 port map( A => n4451, B => n4450, S => n737, Z => n4452);
   U5016 : MUX2_X1 port map( A => n4452, B => n4449, S => n670, Z => n4453);
   U5017 : MUX2_X1 port map( A => REGISTERS_29_24_port, B => 
                           REGISTERS_31_24_port, S => n690, Z => n4454);
   U5018 : MUX2_X1 port map( A => REGISTERS_28_24_port, B => 
                           REGISTERS_30_24_port, S => n690, Z => n4455);
   U5019 : MUX2_X1 port map( A => n4455, B => n4454, S => n737, Z => n4456);
   U5020 : MUX2_X1 port map( A => REGISTERS_25_24_port, B => 
                           REGISTERS_27_24_port, S => n690, Z => n4457);
   U5021 : MUX2_X1 port map( A => REGISTERS_24_24_port, B => 
                           REGISTERS_26_24_port, S => n690, Z => n4458);
   U5022 : MUX2_X1 port map( A => n4458, B => n4457, S => n737, Z => n4459);
   U5023 : MUX2_X1 port map( A => n4459, B => n4456, S => n670, Z => n4460);
   U5024 : MUX2_X1 port map( A => REGISTERS_21_24_port, B => 
                           REGISTERS_23_24_port, S => n690, Z => n4461);
   U5025 : MUX2_X1 port map( A => REGISTERS_20_24_port, B => 
                           REGISTERS_22_24_port, S => n690, Z => n4462);
   U5026 : MUX2_X1 port map( A => n4462, B => n4461, S => n737, Z => n4463);
   U5027 : MUX2_X1 port map( A => REGISTERS_17_24_port, B => 
                           REGISTERS_19_24_port, S => n690, Z => n4464);
   U5028 : MUX2_X1 port map( A => REGISTERS_16_24_port, B => 
                           REGISTERS_18_24_port, S => n690, Z => n4465);
   U5029 : MUX2_X1 port map( A => n4465, B => n4464, S => n737, Z => n4466);
   U5030 : MUX2_X1 port map( A => n4466, B => n4463, S => n670, Z => n4467);
   U5031 : MUX2_X1 port map( A => n4467, B => n4460, S => r3007_A_3_port, Z => 
                           n4468);
   U5032 : MUX2_X1 port map( A => REGISTERS_13_24_port, B => 
                           REGISTERS_15_24_port, S => n689, Z => n4469);
   U5033 : MUX2_X1 port map( A => REGISTERS_12_24_port, B => 
                           REGISTERS_14_24_port, S => n689, Z => n4470);
   U5034 : MUX2_X1 port map( A => n4470, B => n4469, S => n737, Z => n4471);
   U5035 : MUX2_X1 port map( A => REGISTERS_9_24_port, B => 
                           REGISTERS_11_24_port, S => n689, Z => n4472);
   U5036 : MUX2_X1 port map( A => REGISTERS_8_24_port, B => 
                           REGISTERS_10_24_port, S => n689, Z => n4473);
   U5037 : MUX2_X1 port map( A => n4473, B => n4472, S => n736, Z => n4474);
   U5038 : MUX2_X1 port map( A => n4474, B => n4471, S => n670, Z => n4475);
   U5039 : MUX2_X1 port map( A => REGISTERS_5_24_port, B => REGISTERS_7_24_port
                           , S => n689, Z => n4476);
   U5040 : MUX2_X1 port map( A => REGISTERS_4_24_port, B => REGISTERS_6_24_port
                           , S => n689, Z => n4477);
   U5041 : MUX2_X1 port map( A => n4477, B => n4476, S => n736, Z => n4478);
   U5042 : MUX2_X1 port map( A => REGISTERS_1_24_port, B => REGISTERS_3_24_port
                           , S => n689, Z => n4479);
   U5043 : MUX2_X1 port map( A => REGISTERS_0_24_port, B => REGISTERS_2_24_port
                           , S => n689, Z => n4480);
   U5044 : MUX2_X1 port map( A => n4480, B => n4479, S => n736, Z => n4481);
   U5045 : MUX2_X1 port map( A => n4481, B => n4478, S => n670, Z => n4482);
   U5046 : MUX2_X1 port map( A => n4482, B => n4475, S => r3007_A_3_port, Z => 
                           n4483);
   U5047 : MUX2_X1 port map( A => n4483, B => n4468, S => r3007_A_4_port, Z => 
                           n4484);
   U5048 : MUX2_X1 port map( A => n4484, B => n4453, S => ADD_RD1_5_port, Z => 
                           N4396);
   U5049 : MUX2_X1 port map( A => REGISTERS_37_25_port, B => 
                           REGISTERS_39_25_port, S => n689, Z => n4485);
   U5050 : MUX2_X1 port map( A => REGISTERS_36_25_port, B => 
                           REGISTERS_38_25_port, S => n689, Z => n4486);
   U5051 : MUX2_X1 port map( A => n4486, B => n4485, S => n736, Z => n4487);
   U5052 : MUX2_X1 port map( A => REGISTERS_33_25_port, B => 
                           REGISTERS_35_25_port, S => n689, Z => n4488);
   U5053 : MUX2_X1 port map( A => REGISTERS_32_25_port, B => 
                           REGISTERS_34_25_port, S => n689, Z => n4489);
   U5054 : MUX2_X1 port map( A => n4489, B => n4488, S => n736, Z => n4490);
   U5055 : MUX2_X1 port map( A => n4490, B => n4487, S => n670, Z => n4491);
   U5056 : MUX2_X1 port map( A => REGISTERS_29_25_port, B => 
                           REGISTERS_31_25_port, S => n689, Z => n4492);
   U5057 : MUX2_X1 port map( A => REGISTERS_28_25_port, B => 
                           REGISTERS_30_25_port, S => n689, Z => n4493);
   U5058 : MUX2_X1 port map( A => n4493, B => n4492, S => n736, Z => n4494);
   U5059 : MUX2_X1 port map( A => REGISTERS_25_25_port, B => 
                           REGISTERS_27_25_port, S => n689, Z => n4495_port);
   U5060 : MUX2_X1 port map( A => REGISTERS_24_25_port, B => 
                           REGISTERS_26_25_port, S => n688, Z => n4496_port);
   U5061 : MUX2_X1 port map( A => n4496_port, B => n4495_port, S => n736, Z => 
                           n4497_port);
   U5062 : MUX2_X1 port map( A => n4497_port, B => n4494, S => n670, Z => 
                           n4498_port);
   U5063 : MUX2_X1 port map( A => REGISTERS_21_25_port, B => 
                           REGISTERS_23_25_port, S => n688, Z => n4499_port);
   U5064 : MUX2_X1 port map( A => REGISTERS_20_25_port, B => 
                           REGISTERS_22_25_port, S => n688, Z => n4500_port);
   U5065 : MUX2_X1 port map( A => n4500_port, B => n4499_port, S => n736, Z => 
                           n4501_port);
   U5066 : MUX2_X1 port map( A => REGISTERS_17_25_port, B => 
                           REGISTERS_19_25_port, S => n688, Z => n4502_port);
   U5067 : MUX2_X1 port map( A => REGISTERS_16_25_port, B => 
                           REGISTERS_18_25_port, S => n688, Z => n4503_port);
   U5068 : MUX2_X1 port map( A => n4503_port, B => n4502_port, S => n736, Z => 
                           n4504_port);
   U5069 : MUX2_X1 port map( A => n4504_port, B => n4501_port, S => n670, Z => 
                           n4505_port);
   U5070 : MUX2_X1 port map( A => n4505_port, B => n4498_port, S => 
                           r3007_A_3_port, Z => n4506_port);
   U5071 : MUX2_X1 port map( A => REGISTERS_13_25_port, B => 
                           REGISTERS_15_25_port, S => n688, Z => n4507_port);
   U5072 : MUX2_X1 port map( A => REGISTERS_12_25_port, B => 
                           REGISTERS_14_25_port, S => n688, Z => n4508_port);
   U5073 : MUX2_X1 port map( A => n4508_port, B => n4507_port, S => n736, Z => 
                           n4509_port);
   U5074 : MUX2_X1 port map( A => REGISTERS_9_25_port, B => 
                           REGISTERS_11_25_port, S => n688, Z => n4510_port);
   U5075 : MUX2_X1 port map( A => REGISTERS_8_25_port, B => 
                           REGISTERS_10_25_port, S => n688, Z => n4511_port);
   U5076 : MUX2_X1 port map( A => n4511_port, B => n4510_port, S => n736, Z => 
                           n4512_port);
   U5077 : MUX2_X1 port map( A => n4512_port, B => n4509_port, S => n670, Z => 
                           n4513_port);
   U5078 : MUX2_X1 port map( A => REGISTERS_5_25_port, B => REGISTERS_7_25_port
                           , S => n688, Z => n4514_port);
   U5079 : MUX2_X1 port map( A => REGISTERS_4_25_port, B => REGISTERS_6_25_port
                           , S => n688, Z => n4515_port);
   U5080 : MUX2_X1 port map( A => n4515_port, B => n4514_port, S => n736, Z => 
                           n4516_port);
   U5081 : MUX2_X1 port map( A => REGISTERS_1_25_port, B => REGISTERS_3_25_port
                           , S => n688, Z => n4517_port);
   U5082 : MUX2_X1 port map( A => REGISTERS_0_25_port, B => REGISTERS_2_25_port
                           , S => n688, Z => n4518_port);
   U5083 : MUX2_X1 port map( A => n4518_port, B => n4517_port, S => n736, Z => 
                           n4519_port);
   U5084 : MUX2_X1 port map( A => n4519_port, B => n4516_port, S => n670, Z => 
                           n4520_port);
   U5085 : MUX2_X1 port map( A => n4520_port, B => n4513_port, S => 
                           r3007_A_3_port, Z => n4521_port);
   U5086 : MUX2_X1 port map( A => n4521_port, B => n4506_port, S => 
                           r3007_A_4_port, Z => n4522_port);
   U5087 : MUX2_X1 port map( A => n4522_port, B => n4491, S => ADD_RD1_5_port, 
                           Z => N4395);
   U5088 : MUX2_X1 port map( A => REGISTERS_37_26_port, B => 
                           REGISTERS_39_26_port, S => n688, Z => n4523_port);
   U5089 : MUX2_X1 port map( A => REGISTERS_36_26_port, B => 
                           REGISTERS_38_26_port, S => n688, Z => n4524_port);
   U5090 : MUX2_X1 port map( A => n4524_port, B => n4523_port, S => n736, Z => 
                           n4525_port);
   U5091 : MUX2_X1 port map( A => REGISTERS_33_26_port, B => 
                           REGISTERS_35_26_port, S => n687, Z => n4526_port);
   U5092 : MUX2_X1 port map( A => REGISTERS_32_26_port, B => 
                           REGISTERS_34_26_port, S => n687, Z => n4527);
   U5093 : MUX2_X1 port map( A => n4527, B => n4526_port, S => n736, Z => n4528
                           );
   U5094 : MUX2_X1 port map( A => n4528, B => n4525_port, S => n670, Z => n4529
                           );
   U5095 : MUX2_X1 port map( A => REGISTERS_29_26_port, B => 
                           REGISTERS_31_26_port, S => n687, Z => n4530);
   U5096 : MUX2_X1 port map( A => REGISTERS_28_26_port, B => 
                           REGISTERS_30_26_port, S => n687, Z => n4531);
   U5097 : MUX2_X1 port map( A => n4531, B => n4530, S => n735, Z => n4532);
   U5098 : MUX2_X1 port map( A => REGISTERS_25_26_port, B => 
                           REGISTERS_27_26_port, S => n687, Z => n4533);
   U5099 : MUX2_X1 port map( A => REGISTERS_24_26_port, B => 
                           REGISTERS_26_26_port, S => n687, Z => n4534);
   U5100 : MUX2_X1 port map( A => n4534, B => n4533, S => n735, Z => n4535);
   U5101 : MUX2_X1 port map( A => n4535, B => n4532, S => n670, Z => n4536);
   U5102 : MUX2_X1 port map( A => REGISTERS_21_26_port, B => 
                           REGISTERS_23_26_port, S => n687, Z => n4537);
   U5103 : MUX2_X1 port map( A => REGISTERS_20_26_port, B => 
                           REGISTERS_22_26_port, S => n687, Z => n4538);
   U5104 : MUX2_X1 port map( A => n4538, B => n4537, S => n735, Z => n4539);
   U5105 : MUX2_X1 port map( A => REGISTERS_17_26_port, B => 
                           REGISTERS_19_26_port, S => n687, Z => n4540);
   U5106 : MUX2_X1 port map( A => REGISTERS_16_26_port, B => 
                           REGISTERS_18_26_port, S => n687, Z => n4541);
   U5107 : MUX2_X1 port map( A => n4541, B => n4540, S => n735, Z => n4542);
   U5108 : MUX2_X1 port map( A => n4542, B => n4539, S => n670, Z => n4543);
   U5109 : MUX2_X1 port map( A => n4543, B => n4536, S => r3007_A_3_port, Z => 
                           n4544);
   U5110 : MUX2_X1 port map( A => REGISTERS_13_26_port, B => 
                           REGISTERS_15_26_port, S => n687, Z => n4545);
   U5111 : MUX2_X1 port map( A => REGISTERS_12_26_port, B => 
                           REGISTERS_14_26_port, S => n687, Z => n4546);
   U5112 : MUX2_X1 port map( A => n4546, B => n4545, S => n735, Z => n4547);
   U5113 : MUX2_X1 port map( A => REGISTERS_9_26_port, B => 
                           REGISTERS_11_26_port, S => n687, Z => n4548);
   U5114 : MUX2_X1 port map( A => REGISTERS_8_26_port, B => 
                           REGISTERS_10_26_port, S => n687, Z => n4549);
   U5115 : MUX2_X1 port map( A => n4549, B => n4548, S => n735, Z => n4550);
   U5116 : MUX2_X1 port map( A => n4550, B => n4547, S => n669, Z => n4551);
   U5117 : MUX2_X1 port map( A => REGISTERS_5_26_port, B => REGISTERS_7_26_port
                           , S => n687, Z => n4552);
   U5118 : MUX2_X1 port map( A => REGISTERS_4_26_port, B => REGISTERS_6_26_port
                           , S => n686, Z => n4553);
   U5119 : MUX2_X1 port map( A => n4553, B => n4552, S => n735, Z => n4554);
   U5120 : MUX2_X1 port map( A => REGISTERS_1_26_port, B => REGISTERS_3_26_port
                           , S => n686, Z => n4555);
   U5121 : MUX2_X1 port map( A => REGISTERS_0_26_port, B => REGISTERS_2_26_port
                           , S => n686, Z => n4556);
   U5122 : MUX2_X1 port map( A => n4556, B => n4555, S => n735, Z => n4557);
   U5123 : MUX2_X1 port map( A => n4557, B => n4554, S => n669, Z => n4558);
   U5124 : MUX2_X1 port map( A => n4558, B => n4551, S => r3007_A_3_port, Z => 
                           n4559);
   U5125 : MUX2_X1 port map( A => n4559, B => n4544, S => r3007_A_4_port, Z => 
                           n4560);
   U5126 : MUX2_X1 port map( A => n4560, B => n4529, S => ADD_RD1_5_port, Z => 
                           N4394);
   U5127 : MUX2_X1 port map( A => REGISTERS_37_27_port, B => 
                           REGISTERS_39_27_port, S => n686, Z => n4561);
   U5128 : MUX2_X1 port map( A => REGISTERS_36_27_port, B => 
                           REGISTERS_38_27_port, S => n686, Z => n4562);
   U5129 : MUX2_X1 port map( A => n4562, B => n4561, S => n735, Z => n4563);
   U5130 : MUX2_X1 port map( A => REGISTERS_33_27_port, B => 
                           REGISTERS_35_27_port, S => n686, Z => n4564);
   U5131 : MUX2_X1 port map( A => REGISTERS_32_27_port, B => 
                           REGISTERS_34_27_port, S => n686, Z => n4565);
   U5132 : MUX2_X1 port map( A => n4565, B => n4564, S => n735, Z => n4566);
   U5133 : MUX2_X1 port map( A => n4566, B => n4563, S => n669, Z => n4567);
   U5134 : MUX2_X1 port map( A => REGISTERS_29_27_port, B => 
                           REGISTERS_31_27_port, S => n686, Z => n4568);
   U5135 : MUX2_X1 port map( A => REGISTERS_28_27_port, B => 
                           REGISTERS_30_27_port, S => n686, Z => n4569);
   U5136 : MUX2_X1 port map( A => n4569, B => n4568, S => n735, Z => n4570);
   U5137 : MUX2_X1 port map( A => REGISTERS_25_27_port, B => 
                           REGISTERS_27_27_port, S => n686, Z => n4571);
   U5138 : MUX2_X1 port map( A => REGISTERS_24_27_port, B => 
                           REGISTERS_26_27_port, S => n686, Z => n4572);
   U5139 : MUX2_X1 port map( A => n4572, B => n4571, S => n735, Z => n4573);
   U5140 : MUX2_X1 port map( A => n4573, B => n4570, S => n669, Z => n4574);
   U5141 : MUX2_X1 port map( A => REGISTERS_21_27_port, B => 
                           REGISTERS_23_27_port, S => n686, Z => n4575);
   U5142 : MUX2_X1 port map( A => REGISTERS_20_27_port, B => 
                           REGISTERS_22_27_port, S => n686, Z => n4576);
   U5143 : MUX2_X1 port map( A => n4576, B => n4575, S => n735, Z => n4577);
   U5144 : MUX2_X1 port map( A => REGISTERS_17_27_port, B => 
                           REGISTERS_19_27_port, S => n686, Z => n4578);
   U5145 : MUX2_X1 port map( A => REGISTERS_16_27_port, B => 
                           REGISTERS_18_27_port, S => n686, Z => n4579);
   U5146 : MUX2_X1 port map( A => n4579, B => n4578, S => n735, Z => n4580);
   U5147 : MUX2_X1 port map( A => n4580, B => n4577, S => n669, Z => n4581);
   U5148 : MUX2_X1 port map( A => n4581, B => n4574, S => r3007_A_3_port, Z => 
                           n4582);
   U5149 : MUX2_X1 port map( A => REGISTERS_13_27_port, B => 
                           REGISTERS_15_27_port, S => n685, Z => n4583);
   U5150 : MUX2_X1 port map( A => REGISTERS_12_27_port, B => 
                           REGISTERS_14_27_port, S => n685, Z => n4584);
   U5151 : MUX2_X1 port map( A => n4584, B => n4583, S => n735, Z => n4585);
   U5152 : MUX2_X1 port map( A => REGISTERS_9_27_port, B => 
                           REGISTERS_11_27_port, S => n685, Z => n4586);
   U5153 : MUX2_X1 port map( A => REGISTERS_8_27_port, B => 
                           REGISTERS_10_27_port, S => n685, Z => n4587);
   U5154 : MUX2_X1 port map( A => n4587, B => n4586, S => n734, Z => n4588);
   U5155 : MUX2_X1 port map( A => n4588, B => n4585, S => n669, Z => n4589);
   U5156 : MUX2_X1 port map( A => REGISTERS_5_27_port, B => REGISTERS_7_27_port
                           , S => n685, Z => n4590);
   U5157 : MUX2_X1 port map( A => REGISTERS_4_27_port, B => REGISTERS_6_27_port
                           , S => n685, Z => n4591);
   U5158 : MUX2_X1 port map( A => n4591, B => n4590, S => n734, Z => n4592);
   U5159 : MUX2_X1 port map( A => REGISTERS_1_27_port, B => REGISTERS_3_27_port
                           , S => n685, Z => n4593);
   U5160 : MUX2_X1 port map( A => REGISTERS_0_27_port, B => REGISTERS_2_27_port
                           , S => n685, Z => n4594);
   U5161 : MUX2_X1 port map( A => n4594, B => n4593, S => n734, Z => n4595);
   U5162 : MUX2_X1 port map( A => n4595, B => n4592, S => n669, Z => n4596);
   U5163 : MUX2_X1 port map( A => n4596, B => n4589, S => r3007_A_3_port, Z => 
                           n4597);
   U5164 : MUX2_X1 port map( A => n4597, B => n4582, S => r3007_A_4_port, Z => 
                           n4598);
   U5165 : MUX2_X1 port map( A => n4598, B => n4567, S => ADD_RD1_5_port, Z => 
                           N4393);
   U5166 : MUX2_X1 port map( A => REGISTERS_37_28_port, B => 
                           REGISTERS_39_28_port, S => n685, Z => n4599);
   U5167 : MUX2_X1 port map( A => REGISTERS_36_28_port, B => 
                           REGISTERS_38_28_port, S => n685, Z => n4600);
   U5168 : MUX2_X1 port map( A => n4600, B => n4599, S => n734, Z => n4601);
   U5169 : MUX2_X1 port map( A => REGISTERS_33_28_port, B => 
                           REGISTERS_35_28_port, S => n685, Z => n4602);
   U5170 : MUX2_X1 port map( A => REGISTERS_32_28_port, B => 
                           REGISTERS_34_28_port, S => n685, Z => n4603);
   U5171 : MUX2_X1 port map( A => n4603, B => n4602, S => n734, Z => n4604);
   U5172 : MUX2_X1 port map( A => n4604, B => n4601, S => n669, Z => n4605);
   U5173 : MUX2_X1 port map( A => REGISTERS_29_28_port, B => 
                           REGISTERS_31_28_port, S => n685, Z => n4606);
   U5174 : MUX2_X1 port map( A => REGISTERS_28_28_port, B => 
                           REGISTERS_30_28_port, S => n685, Z => n4607);
   U5175 : MUX2_X1 port map( A => n4607, B => n4606, S => n734, Z => n4608);
   U5176 : MUX2_X1 port map( A => REGISTERS_25_28_port, B => 
                           REGISTERS_27_28_port, S => n685, Z => n4609);
   U5177 : MUX2_X1 port map( A => REGISTERS_24_28_port, B => 
                           REGISTERS_26_28_port, S => n684, Z => n4610);
   U5178 : MUX2_X1 port map( A => n4610, B => n4609, S => n734, Z => n4611);
   U5179 : MUX2_X1 port map( A => n4611, B => n4608, S => n669, Z => n4612);
   U5180 : MUX2_X1 port map( A => REGISTERS_21_28_port, B => 
                           REGISTERS_23_28_port, S => n684, Z => n4613);
   U5181 : MUX2_X1 port map( A => REGISTERS_20_28_port, B => 
                           REGISTERS_22_28_port, S => n684, Z => n4614);
   U5182 : MUX2_X1 port map( A => n4614, B => n4613, S => n734, Z => n4615);
   U5183 : MUX2_X1 port map( A => REGISTERS_17_28_port, B => 
                           REGISTERS_19_28_port, S => n684, Z => n4616);
   U5184 : MUX2_X1 port map( A => REGISTERS_16_28_port, B => 
                           REGISTERS_18_28_port, S => n684, Z => n4617);
   U5185 : MUX2_X1 port map( A => n4617, B => n4616, S => n734, Z => n4618);
   U5186 : MUX2_X1 port map( A => n4618, B => n4615, S => n669, Z => n4619);
   U5187 : MUX2_X1 port map( A => n4619, B => n4612, S => r3007_A_3_port, Z => 
                           n4620);
   U5188 : MUX2_X1 port map( A => REGISTERS_13_28_port, B => 
                           REGISTERS_15_28_port, S => n684, Z => n4621);
   U5189 : MUX2_X1 port map( A => REGISTERS_12_28_port, B => 
                           REGISTERS_14_28_port, S => n684, Z => n4622);
   U5190 : MUX2_X1 port map( A => n4622, B => n4621, S => n734, Z => n4623);
   U5191 : MUX2_X1 port map( A => REGISTERS_9_28_port, B => 
                           REGISTERS_11_28_port, S => n684, Z => n4624);
   U5192 : MUX2_X1 port map( A => REGISTERS_8_28_port, B => 
                           REGISTERS_10_28_port, S => n684, Z => n4625);
   U5193 : MUX2_X1 port map( A => n4625, B => n4624, S => n734, Z => n4626);
   U5194 : MUX2_X1 port map( A => n4626, B => n4623, S => n669, Z => n4627);
   U5195 : MUX2_X1 port map( A => REGISTERS_5_28_port, B => REGISTERS_7_28_port
                           , S => n684, Z => n4628);
   U5196 : MUX2_X1 port map( A => REGISTERS_4_28_port, B => REGISTERS_6_28_port
                           , S => n684, Z => n4629);
   U5197 : MUX2_X1 port map( A => n4629, B => n4628, S => n734, Z => n4630);
   U5198 : MUX2_X1 port map( A => REGISTERS_1_28_port, B => REGISTERS_3_28_port
                           , S => n684, Z => n4631);
   U5199 : MUX2_X1 port map( A => REGISTERS_0_28_port, B => REGISTERS_2_28_port
                           , S => n684, Z => n4632);
   U5200 : MUX2_X1 port map( A => n4632, B => n4631, S => n734, Z => n4633);
   U5201 : MUX2_X1 port map( A => n4633, B => n4630, S => n669, Z => n4634);
   U5202 : MUX2_X1 port map( A => n4634, B => n4627, S => r3007_A_3_port, Z => 
                           n4635);
   U5203 : MUX2_X1 port map( A => n4635, B => n4620, S => r3007_A_4_port, Z => 
                           n4636);
   U5204 : MUX2_X1 port map( A => n4636, B => n4605, S => ADD_RD1_5_port, Z => 
                           N4392);
   U5205 : MUX2_X1 port map( A => REGISTERS_37_29_port, B => 
                           REGISTERS_39_29_port, S => n684, Z => n4637);
   U5206 : MUX2_X1 port map( A => REGISTERS_36_29_port, B => 
                           REGISTERS_38_29_port, S => n684, Z => n4638);
   U5207 : MUX2_X1 port map( A => n4638, B => n4637, S => n734, Z => n4639);
   U5208 : MUX2_X1 port map( A => REGISTERS_33_29_port, B => 
                           REGISTERS_35_29_port, S => n683, Z => n4640);
   U5209 : MUX2_X1 port map( A => REGISTERS_32_29_port, B => 
                           REGISTERS_34_29_port, S => n683, Z => n4641);
   U5210 : MUX2_X1 port map( A => n4641, B => n4640, S => n734, Z => n4642);
   U5211 : MUX2_X1 port map( A => n4642, B => n4639, S => n669, Z => n4643);
   U5212 : MUX2_X1 port map( A => REGISTERS_29_29_port, B => 
                           REGISTERS_31_29_port, S => n683, Z => n4644);
   U5213 : MUX2_X1 port map( A => REGISTERS_28_29_port, B => 
                           REGISTERS_30_29_port, S => n683, Z => n4645);
   U5214 : MUX2_X1 port map( A => n4645, B => n4644, S => n733, Z => n4646);
   U5215 : MUX2_X1 port map( A => REGISTERS_25_29_port, B => 
                           REGISTERS_27_29_port, S => n683, Z => n4647);
   U5216 : MUX2_X1 port map( A => REGISTERS_24_29_port, B => 
                           REGISTERS_26_29_port, S => n683, Z => n4648);
   U5217 : MUX2_X1 port map( A => n4648, B => n4647, S => n733, Z => n4649);
   U5218 : MUX2_X1 port map( A => n4649, B => n4646, S => n669, Z => n4650);
   U5219 : MUX2_X1 port map( A => REGISTERS_21_29_port, B => 
                           REGISTERS_23_29_port, S => n683, Z => n4651);
   U5220 : MUX2_X1 port map( A => REGISTERS_20_29_port, B => 
                           REGISTERS_22_29_port, S => n683, Z => n4652);
   U5221 : MUX2_X1 port map( A => n4652, B => n4651, S => n733, Z => n4653);
   U5222 : MUX2_X1 port map( A => REGISTERS_17_29_port, B => 
                           REGISTERS_19_29_port, S => n683, Z => n4654);
   U5223 : MUX2_X1 port map( A => REGISTERS_16_29_port, B => 
                           REGISTERS_18_29_port, S => n683, Z => n4655);
   U5224 : MUX2_X1 port map( A => n4655, B => n4654, S => n733, Z => n4656);
   U5225 : MUX2_X1 port map( A => n4656, B => n4653, S => n668, Z => n4657);
   U5226 : MUX2_X1 port map( A => n4657, B => n4650, S => r3007_A_3_port, Z => 
                           n4658);
   U5227 : MUX2_X1 port map( A => REGISTERS_13_29_port, B => 
                           REGISTERS_15_29_port, S => n683, Z => n4659);
   U5228 : MUX2_X1 port map( A => REGISTERS_12_29_port, B => 
                           REGISTERS_14_29_port, S => n683, Z => n4660);
   U5229 : MUX2_X1 port map( A => n4660, B => n4659, S => n733, Z => n4661);
   U5230 : MUX2_X1 port map( A => REGISTERS_9_29_port, B => 
                           REGISTERS_11_29_port, S => n683, Z => n4662);
   U5231 : MUX2_X1 port map( A => REGISTERS_8_29_port, B => 
                           REGISTERS_10_29_port, S => n683, Z => n4663);
   U5232 : MUX2_X1 port map( A => n4663, B => n4662, S => n733, Z => n4664);
   U5233 : MUX2_X1 port map( A => n4664, B => n4661, S => n668, Z => n4665);
   U5234 : MUX2_X1 port map( A => REGISTERS_5_29_port, B => REGISTERS_7_29_port
                           , S => n683, Z => n4666);
   U5235 : MUX2_X1 port map( A => REGISTERS_4_29_port, B => REGISTERS_6_29_port
                           , S => n682, Z => n4667);
   U5236 : MUX2_X1 port map( A => n4667, B => n4666, S => n733, Z => n4668);
   U5237 : MUX2_X1 port map( A => REGISTERS_1_29_port, B => REGISTERS_3_29_port
                           , S => n682, Z => n4669);
   U5238 : MUX2_X1 port map( A => REGISTERS_0_29_port, B => REGISTERS_2_29_port
                           , S => n682, Z => n4670);
   U5239 : MUX2_X1 port map( A => n4670, B => n4669, S => n733, Z => n4671);
   U5240 : MUX2_X1 port map( A => n4671, B => n4668, S => n668, Z => n4672);
   U5241 : MUX2_X1 port map( A => n4672, B => n4665, S => r3007_A_3_port, Z => 
                           n4673);
   U5242 : MUX2_X1 port map( A => n4673, B => n4658, S => r3007_A_4_port, Z => 
                           n4674);
   U5243 : MUX2_X1 port map( A => n4674, B => n4643, S => ADD_RD1_5_port, Z => 
                           N4391);
   U5244 : MUX2_X1 port map( A => REGISTERS_37_30_port, B => 
                           REGISTERS_39_30_port, S => n682, Z => n4675);
   U5245 : MUX2_X1 port map( A => REGISTERS_36_30_port, B => 
                           REGISTERS_38_30_port, S => n682, Z => n4676);
   U5246 : MUX2_X1 port map( A => n4676, B => n4675, S => n733, Z => n4677);
   U5247 : MUX2_X1 port map( A => REGISTERS_33_30_port, B => 
                           REGISTERS_35_30_port, S => n682, Z => n4678);
   U5248 : MUX2_X1 port map( A => REGISTERS_32_30_port, B => 
                           REGISTERS_34_30_port, S => n682, Z => n4679);
   U5249 : MUX2_X1 port map( A => n4679, B => n4678, S => n733, Z => n4680);
   U5250 : MUX2_X1 port map( A => n4680, B => n4677, S => n668, Z => n4681);
   U5251 : MUX2_X1 port map( A => REGISTERS_29_30_port, B => 
                           REGISTERS_31_30_port, S => n682, Z => n4682);
   U5252 : MUX2_X1 port map( A => REGISTERS_28_30_port, B => 
                           REGISTERS_30_30_port, S => n682, Z => n4683);
   U5253 : MUX2_X1 port map( A => n4683, B => n4682, S => n733, Z => n4684);
   U5254 : MUX2_X1 port map( A => REGISTERS_25_30_port, B => 
                           REGISTERS_27_30_port, S => n682, Z => n4685);
   U5255 : MUX2_X1 port map( A => REGISTERS_24_30_port, B => 
                           REGISTERS_26_30_port, S => n682, Z => n4686);
   U5256 : MUX2_X1 port map( A => n4686, B => n4685, S => n733, Z => n4687);
   U5257 : MUX2_X1 port map( A => n4687, B => n4684, S => n668, Z => n4688);
   U5258 : MUX2_X1 port map( A => REGISTERS_21_30_port, B => 
                           REGISTERS_23_30_port, S => n682, Z => n4689);
   U5259 : MUX2_X1 port map( A => REGISTERS_20_30_port, B => 
                           REGISTERS_22_30_port, S => n682, Z => n4690);
   U5260 : MUX2_X1 port map( A => n4690, B => n4689, S => n733, Z => n4691);
   U5261 : MUX2_X1 port map( A => REGISTERS_17_30_port, B => 
                           REGISTERS_19_30_port, S => n682, Z => n4692);
   U5262 : MUX2_X1 port map( A => REGISTERS_16_30_port, B => 
                           REGISTERS_18_30_port, S => n682, Z => n4693);
   U5263 : MUX2_X1 port map( A => n4693, B => n4692, S => n733, Z => n4694);
   U5264 : MUX2_X1 port map( A => n4694, B => n4691, S => n668, Z => n4695);
   U5265 : MUX2_X1 port map( A => n4695, B => n4688, S => r3007_A_3_port, Z => 
                           n4696);
   U5266 : MUX2_X1 port map( A => REGISTERS_13_30_port, B => 
                           REGISTERS_15_30_port, S => n681, Z => n4697);
   U5267 : MUX2_X1 port map( A => REGISTERS_12_30_port, B => 
                           REGISTERS_14_30_port, S => n681, Z => n4698);
   U5268 : MUX2_X1 port map( A => n4698, B => n4697, S => n733, Z => n4699);
   U5269 : MUX2_X1 port map( A => REGISTERS_9_30_port, B => 
                           REGISTERS_11_30_port, S => n681, Z => n4700);
   U5270 : MUX2_X1 port map( A => REGISTERS_8_30_port, B => 
                           REGISTERS_10_30_port, S => n681, Z => n4701);
   U5271 : MUX2_X1 port map( A => n4701, B => n4700, S => n732, Z => n4702);
   U5272 : MUX2_X1 port map( A => n4702, B => n4699, S => n668, Z => n4703);
   U5273 : MUX2_X1 port map( A => REGISTERS_5_30_port, B => REGISTERS_7_30_port
                           , S => n681, Z => n4704);
   U5274 : MUX2_X1 port map( A => REGISTERS_4_30_port, B => REGISTERS_6_30_port
                           , S => n681, Z => n4705);
   U5275 : MUX2_X1 port map( A => n4705, B => n4704, S => n732, Z => n4706);
   U5276 : MUX2_X1 port map( A => REGISTERS_1_30_port, B => REGISTERS_3_30_port
                           , S => n681, Z => n4707);
   U5277 : MUX2_X1 port map( A => REGISTERS_0_30_port, B => REGISTERS_2_30_port
                           , S => n681, Z => n4708);
   U5278 : MUX2_X1 port map( A => n4708, B => n4707, S => n732, Z => n4709);
   U5279 : MUX2_X1 port map( A => n4709, B => n4706, S => n668, Z => n4710);
   U5280 : MUX2_X1 port map( A => n4710, B => n4703, S => r3007_A_3_port, Z => 
                           n4711);
   U5281 : MUX2_X1 port map( A => n4711, B => n4696, S => r3007_A_4_port, Z => 
                           n4712);
   U5282 : MUX2_X1 port map( A => n4712, B => n4681, S => ADD_RD1_5_port, Z => 
                           N4390);
   U5283 : MUX2_X1 port map( A => REGISTERS_37_31_port, B => 
                           REGISTERS_39_31_port, S => n681, Z => n4713);
   U5284 : MUX2_X1 port map( A => REGISTERS_36_31_port, B => 
                           REGISTERS_38_31_port, S => n681, Z => n4714);
   U5285 : MUX2_X1 port map( A => n4714, B => n4713, S => n732, Z => n4715);
   U5286 : MUX2_X1 port map( A => REGISTERS_33_31_port, B => 
                           REGISTERS_35_31_port, S => n681, Z => n4716);
   U5287 : MUX2_X1 port map( A => REGISTERS_32_31_port, B => 
                           REGISTERS_34_31_port, S => n681, Z => n4717);
   U5288 : MUX2_X1 port map( A => n4717, B => n4716, S => n732, Z => n4718);
   U5289 : MUX2_X1 port map( A => n4718, B => n4715, S => n668, Z => n4719);
   U5290 : MUX2_X1 port map( A => REGISTERS_29_31_port, B => 
                           REGISTERS_31_31_port, S => n681, Z => n4720);
   U5291 : MUX2_X1 port map( A => REGISTERS_28_31_port, B => 
                           REGISTERS_30_31_port, S => n681, Z => n4721);
   U5292 : MUX2_X1 port map( A => n4721, B => n4720, S => n732, Z => n4722);
   U5293 : MUX2_X1 port map( A => REGISTERS_25_31_port, B => 
                           REGISTERS_27_31_port, S => n681, Z => n4723);
   U5294 : MUX2_X1 port map( A => REGISTERS_24_31_port, B => 
                           REGISTERS_26_31_port, S => n680, Z => n4724);
   U5295 : MUX2_X1 port map( A => n4724, B => n4723, S => n732, Z => n4725);
   U5296 : MUX2_X1 port map( A => n4725, B => n4722, S => n668, Z => n4726);
   U5297 : MUX2_X1 port map( A => REGISTERS_21_31_port, B => 
                           REGISTERS_23_31_port, S => n680, Z => n4727);
   U5298 : MUX2_X1 port map( A => REGISTERS_20_31_port, B => 
                           REGISTERS_22_31_port, S => n680, Z => n4728);
   U5299 : MUX2_X1 port map( A => n4728, B => n4727, S => n732, Z => n4729);
   U5300 : MUX2_X1 port map( A => REGISTERS_17_31_port, B => 
                           REGISTERS_19_31_port, S => n680, Z => n4730);
   U5301 : MUX2_X1 port map( A => REGISTERS_16_31_port, B => 
                           REGISTERS_18_31_port, S => n680, Z => n4731);
   U5302 : MUX2_X1 port map( A => n4731, B => n4730, S => n732, Z => n4732);
   U5303 : MUX2_X1 port map( A => n4732, B => n4729, S => n668, Z => n4733);
   U5304 : MUX2_X1 port map( A => n4733, B => n4726, S => r3007_A_3_port, Z => 
                           n4734);
   U5305 : MUX2_X1 port map( A => REGISTERS_13_31_port, B => 
                           REGISTERS_15_31_port, S => n680, Z => n4735);
   U5306 : MUX2_X1 port map( A => REGISTERS_12_31_port, B => 
                           REGISTERS_14_31_port, S => n680, Z => n4736);
   U5307 : MUX2_X1 port map( A => n4736, B => n4735, S => n732, Z => n4737);
   U5308 : MUX2_X1 port map( A => REGISTERS_9_31_port, B => 
                           REGISTERS_11_31_port, S => n680, Z => n4738);
   U5309 : MUX2_X1 port map( A => REGISTERS_8_31_port, B => 
                           REGISTERS_10_31_port, S => n680, Z => n4739);
   U5310 : MUX2_X1 port map( A => n4739, B => n4738, S => n732, Z => n4740);
   U5311 : MUX2_X1 port map( A => n4740, B => n4737, S => n668, Z => n4741);
   U5312 : MUX2_X1 port map( A => REGISTERS_5_31_port, B => REGISTERS_7_31_port
                           , S => n680, Z => n4742);
   U5313 : MUX2_X1 port map( A => REGISTERS_4_31_port, B => REGISTERS_6_31_port
                           , S => n680, Z => n4743);
   U5314 : MUX2_X1 port map( A => n4743, B => n4742, S => n732, Z => n4744);
   U5315 : MUX2_X1 port map( A => REGISTERS_1_31_port, B => REGISTERS_3_31_port
                           , S => n680, Z => n4745);
   U5316 : MUX2_X1 port map( A => REGISTERS_0_31_port, B => REGISTERS_2_31_port
                           , S => n680, Z => n4746);
   U5317 : MUX2_X1 port map( A => n4746, B => n4745, S => n732, Z => n4747);
   U5318 : MUX2_X1 port map( A => n4747, B => n4744, S => n668, Z => n4748);
   U5319 : MUX2_X1 port map( A => n4748, B => n4741, S => r3007_A_3_port, Z => 
                           n4749);
   U5320 : MUX2_X1 port map( A => n4749, B => n4734, S => r3007_A_4_port, Z => 
                           n4750);
   U5321 : MUX2_X1 port map( A => n4750, B => n4719, S => ADD_RD1_5_port, Z => 
                           N4389);
   U5322 : INV_X1 port map( A => n4751, ZN => n16456);
   U5323 : AOI222_X1 port map( A1 => MEM_OUT_31_port, A2 => n4752, B1 => N5281,
                           B2 => n169, C1 => N12236, C2 => n166, ZN => n4751);
   U5324 : INV_X1 port map( A => n4753, ZN => n16457);
   U5325 : AOI222_X1 port map( A1 => MEM_OUT_30_port, A2 => n4752, B1 => N5280,
                           B2 => n169, C1 => N12235, C2 => n166, ZN => n4753);
   U5326 : INV_X1 port map( A => n4754, ZN => n16458);
   U5327 : AOI222_X1 port map( A1 => MEM_OUT_29_port, A2 => n4752, B1 => N5279,
                           B2 => n169, C1 => N12234, C2 => n166, ZN => n4754);
   U5328 : INV_X1 port map( A => n4755, ZN => n16459);
   U5329 : AOI222_X1 port map( A1 => MEM_OUT_28_port, A2 => n4752, B1 => N5278,
                           B2 => n169, C1 => N12233, C2 => n166, ZN => n4755);
   U5330 : INV_X1 port map( A => n4756, ZN => n16460);
   U5331 : AOI222_X1 port map( A1 => MEM_OUT_27_port, A2 => n4752, B1 => N5277,
                           B2 => n169, C1 => N12232, C2 => n166, ZN => n4756);
   U5332 : INV_X1 port map( A => n4757, ZN => n16461);
   U5333 : AOI222_X1 port map( A1 => MEM_OUT_26_port, A2 => n4752, B1 => N5276,
                           B2 => n169, C1 => N12231, C2 => n166, ZN => n4757);
   U5334 : INV_X1 port map( A => n4758, ZN => n16462);
   U5335 : AOI222_X1 port map( A1 => MEM_OUT_25_port, A2 => n4752, B1 => N5275,
                           B2 => n169, C1 => N12230, C2 => n166, ZN => n4758);
   U5336 : INV_X1 port map( A => n4759, ZN => n16463);
   U5337 : AOI222_X1 port map( A1 => MEM_OUT_24_port, A2 => n4752, B1 => N5274,
                           B2 => n169, C1 => N12229, C2 => n166, ZN => n4759);
   U5338 : INV_X1 port map( A => n4760, ZN => n16464);
   U5339 : AOI222_X1 port map( A1 => MEM_OUT_23_port, A2 => n4752, B1 => N5273,
                           B2 => n169, C1 => N12228, C2 => n166, ZN => n4760);
   U5340 : INV_X1 port map( A => n4761, ZN => n16465);
   U5341 : AOI222_X1 port map( A1 => MEM_OUT_22_port, A2 => n4752, B1 => N5272,
                           B2 => n169, C1 => N12227, C2 => n166, ZN => n4761);
   U5342 : INV_X1 port map( A => n4762, ZN => n16466);
   U5343 : AOI222_X1 port map( A1 => MEM_OUT_21_port, A2 => n4752, B1 => N5271,
                           B2 => n169, C1 => N12226, C2 => n166, ZN => n4762);
   U5344 : INV_X1 port map( A => n4763, ZN => n16467);
   U5345 : AOI222_X1 port map( A1 => MEM_OUT_20_port, A2 => n4752, B1 => N5270,
                           B2 => n169, C1 => N12225, C2 => n166, ZN => n4763);
   U5346 : INV_X1 port map( A => n4764, ZN => n16468);
   U5347 : AOI222_X1 port map( A1 => MEM_OUT_19_port, A2 => n4752, B1 => N5269,
                           B2 => n169, C1 => N12224, C2 => n166, ZN => n4764);
   U5348 : INV_X1 port map( A => n4765, ZN => n16469);
   U5349 : AOI222_X1 port map( A1 => MEM_OUT_18_port, A2 => n4752, B1 => N5268,
                           B2 => n169, C1 => N12223, C2 => n166, ZN => n4765);
   U5350 : INV_X1 port map( A => n4766, ZN => n16470);
   U5351 : AOI222_X1 port map( A1 => MEM_OUT_17_port, A2 => n4752, B1 => N5267,
                           B2 => n169, C1 => N12222, C2 => n166, ZN => n4766);
   U5352 : INV_X1 port map( A => n4767, ZN => n16471);
   U5353 : AOI222_X1 port map( A1 => MEM_OUT_16_port, A2 => n4752, B1 => N5266,
                           B2 => n169, C1 => N12221, C2 => n166, ZN => n4767);
   U5354 : INV_X1 port map( A => n4768, ZN => n16472);
   U5355 : AOI222_X1 port map( A1 => MEM_OUT_15_port, A2 => n4752, B1 => N5265,
                           B2 => n169, C1 => N12220, C2 => n166, ZN => n4768);
   U5356 : INV_X1 port map( A => n4769, ZN => n16473);
   U5357 : AOI222_X1 port map( A1 => MEM_OUT_14_port, A2 => n4752, B1 => N5264,
                           B2 => n169, C1 => N12219, C2 => n166, ZN => n4769);
   U5358 : INV_X1 port map( A => n4770, ZN => n16474);
   U5359 : AOI222_X1 port map( A1 => MEM_OUT_13_port, A2 => n4752, B1 => N5263,
                           B2 => n169, C1 => N12218, C2 => n166, ZN => n4770);
   U5360 : INV_X1 port map( A => n4771, ZN => n16475);
   U5361 : AOI222_X1 port map( A1 => MEM_OUT_12_port, A2 => n4752, B1 => N5262,
                           B2 => n169, C1 => N12217, C2 => n166, ZN => n4771);
   U5362 : INV_X1 port map( A => n4772, ZN => n16476);
   U5363 : AOI222_X1 port map( A1 => MEM_OUT_11_port, A2 => n4752, B1 => N5261,
                           B2 => n169, C1 => N12216, C2 => n166, ZN => n4772);
   U5364 : INV_X1 port map( A => n4773, ZN => n16477);
   U5365 : AOI222_X1 port map( A1 => MEM_OUT_10_port, A2 => n4752, B1 => N5260,
                           B2 => n169, C1 => N12215, C2 => n166, ZN => n4773);
   U5366 : INV_X1 port map( A => n4774, ZN => n16478);
   U5367 : AOI222_X1 port map( A1 => MEM_OUT_9_port, A2 => n4752, B1 => N5259, 
                           B2 => n169, C1 => N12214, C2 => n166, ZN => n4774);
   U5368 : INV_X1 port map( A => n4775, ZN => n16479);
   U5369 : AOI222_X1 port map( A1 => MEM_OUT_8_port, A2 => n4752, B1 => N5258, 
                           B2 => n169, C1 => N12213, C2 => n166, ZN => n4775);
   U5370 : INV_X1 port map( A => n4776, ZN => n16480);
   U5371 : AOI222_X1 port map( A1 => MEM_OUT_7_port, A2 => n4752, B1 => N5257, 
                           B2 => n169, C1 => N12212, C2 => n166, ZN => n4776);
   U5372 : INV_X1 port map( A => n4777, ZN => n16481);
   U5373 : AOI222_X1 port map( A1 => MEM_OUT_6_port, A2 => n4752, B1 => N5256, 
                           B2 => n169, C1 => N12211, C2 => n166, ZN => n4777);
   U5374 : INV_X1 port map( A => n4778, ZN => n16482);
   U5375 : AOI222_X1 port map( A1 => MEM_OUT_5_port, A2 => n4752, B1 => N5255, 
                           B2 => n169, C1 => N12210, C2 => n166, ZN => n4778);
   U5376 : INV_X1 port map( A => n4779, ZN => n16483);
   U5377 : AOI222_X1 port map( A1 => MEM_OUT_4_port, A2 => n4752, B1 => N5254, 
                           B2 => n169, C1 => N12209, C2 => n166, ZN => n4779);
   U5378 : INV_X1 port map( A => n4780, ZN => n16484);
   U5379 : AOI222_X1 port map( A1 => MEM_OUT_3_port, A2 => n4752, B1 => N5253, 
                           B2 => n169, C1 => N12208, C2 => n166, ZN => n4780);
   U5380 : INV_X1 port map( A => n4781, ZN => n16485);
   U5381 : AOI222_X1 port map( A1 => MEM_OUT_2_port, A2 => n4752, B1 => N5252, 
                           B2 => n169, C1 => N12207, C2 => n166, ZN => n4781);
   U5382 : INV_X1 port map( A => n4782, ZN => n16486);
   U5383 : AOI222_X1 port map( A1 => MEM_OUT_1_port, A2 => n4752, B1 => N5251, 
                           B2 => n169, C1 => N12206, C2 => n166, ZN => n4782);
   U5384 : INV_X1 port map( A => n4783, ZN => n16487);
   U5385 : AOI222_X1 port map( A1 => MEM_OUT_0_port, A2 => n4752, B1 => N5250, 
                           B2 => n169, C1 => N12205, C2 => n166, ZN => n4783);
   U5386 : OAI22_X1 port map( A1 => n4786, A2 => n4787, B1 => n4788, B2 => n116
                           , ZN => n13192);
   U5387 : OAI21_X1 port map( B1 => n11790, B2 => n4789, A => n4790, ZN => 
                           n13191);
   U5388 : AOI22_X1 port map( A1 => N13862, A2 => n4791, B1 => N12300, B2 => 
                           n305, ZN => n4790);
   U5389 : OAI21_X1 port map( B1 => n11863, B2 => n4789, A => n4793, ZN => 
                           n13190);
   U5390 : AOI22_X1 port map( A1 => N13831, A2 => n4791, B1 => N12269, B2 => 
                           n305, ZN => n4793);
   U5391 : OAI21_X1 port map( B1 => n11862, B2 => n4789, A => n4794, ZN => 
                           n13189);
   U5392 : AOI22_X1 port map( A1 => N13832, A2 => n4791, B1 => N12270, B2 => 
                           n305, ZN => n4794);
   U5393 : OAI211_X1 port map( C1 => n4795, C2 => n4796, A => n4797, B => n4798
                           , ZN => n13188);
   U5394 : AOI22_X1 port map( A1 => N13833, A2 => n4799, B1 => n4800, B2 => 
                           CWP_2_port, ZN => n4798);
   U5395 : INV_X1 port map( A => n4801, ZN => n4796);
   U5396 : NOR2_X1 port map( A1 => n4802, A2 => N12271, ZN => n4795);
   U5397 : NAND3_X1 port map( A1 => n4803, A2 => n4797, A3 => n4804, ZN => 
                           n13187);
   U5398 : AOI22_X1 port map( A1 => N13834, A2 => n4799, B1 => n4800, B2 => 
                           CWP_3_port, ZN => n4804);
   U5399 : NAND3_X1 port map( A1 => n4801, A2 => n4805, A3 => N12272, ZN => 
                           n4803);
   U5400 : NAND3_X1 port map( A1 => n4806, A2 => n4797, A3 => n4807, ZN => 
                           n13186);
   U5401 : AOI22_X1 port map( A1 => N13835, A2 => n4799, B1 => n4800, B2 => 
                           CWP_4_port, ZN => n4807);
   U5402 : AOI21_X1 port map( B1 => n4808, B2 => n4809, A => n4800, ZN => n4799
                           );
   U5403 : NAND3_X1 port map( A1 => n300, A2 => n4810, A3 => n4789, ZN => n4797
                           );
   U5404 : NAND3_X1 port map( A1 => n4801, A2 => n4805, A3 => N12273, ZN => 
                           n4806);
   U5405 : INV_X1 port map( A => n4802, ZN => n4805);
   U5406 : NOR3_X1 port map( A1 => n4811, A2 => n4812, A3 => n4800, ZN => n4801
                           );
   U5407 : OAI21_X1 port map( B1 => n11842, B2 => n4789, A => n4813, ZN => 
                           n13185);
   U5408 : AOI22_X1 port map( A1 => N13836, A2 => n4791, B1 => N12274, B2 => 
                           n305, ZN => n4813);
   U5409 : OAI21_X1 port map( B1 => n11841, B2 => n4789, A => n4814, ZN => 
                           n13184);
   U5410 : AOI22_X1 port map( A1 => N13837, A2 => n4791, B1 => N12275, B2 => 
                           n305, ZN => n4814);
   U5411 : OAI21_X1 port map( B1 => n11840, B2 => n4789, A => n4815, ZN => 
                           n13183);
   U5412 : AOI22_X1 port map( A1 => N13838, A2 => n4791, B1 => N12276, B2 => 
                           n305, ZN => n4815);
   U5413 : OAI21_X1 port map( B1 => n11839, B2 => n4789, A => n4816, ZN => 
                           n13182);
   U5414 : AOI22_X1 port map( A1 => N13839, A2 => n4791, B1 => N12277, B2 => 
                           n305, ZN => n4816);
   U5415 : OAI21_X1 port map( B1 => n11838, B2 => n4789, A => n4817, ZN => 
                           n13181);
   U5416 : AOI22_X1 port map( A1 => N13840, A2 => n4791, B1 => N12278, B2 => 
                           n305, ZN => n4817);
   U5417 : OAI21_X1 port map( B1 => n11837, B2 => n4789, A => n4818, ZN => 
                           n13180);
   U5418 : AOI22_X1 port map( A1 => N13841, A2 => n4791, B1 => N12279, B2 => 
                           n305, ZN => n4818);
   U5419 : OAI21_X1 port map( B1 => n11836, B2 => n4789, A => n4819, ZN => 
                           n13179);
   U5420 : AOI22_X1 port map( A1 => N13842, A2 => n4791, B1 => N12280, B2 => 
                           n305, ZN => n4819);
   U5421 : OAI21_X1 port map( B1 => n11835, B2 => n4789, A => n4820, ZN => 
                           n13178);
   U5422 : AOI22_X1 port map( A1 => N13843, A2 => n4791, B1 => N12281, B2 => 
                           n305, ZN => n4820);
   U5423 : OAI21_X1 port map( B1 => n11834, B2 => n4789, A => n4821, ZN => 
                           n13177);
   U5424 : AOI22_X1 port map( A1 => N13844, A2 => n4791, B1 => N12282, B2 => 
                           n305, ZN => n4821);
   U5425 : OAI21_X1 port map( B1 => n11833, B2 => n4789, A => n4822, ZN => 
                           n13176);
   U5426 : AOI22_X1 port map( A1 => N13845, A2 => n4791, B1 => N12283, B2 => 
                           n305, ZN => n4822);
   U5427 : OAI21_X1 port map( B1 => n11832, B2 => n4789, A => n4823, ZN => 
                           n13175);
   U5428 : AOI22_X1 port map( A1 => N13846, A2 => n4791, B1 => N12284, B2 => 
                           n305, ZN => n4823);
   U5429 : OAI21_X1 port map( B1 => n11831, B2 => n4789, A => n4824, ZN => 
                           n13174);
   U5430 : AOI22_X1 port map( A1 => N13847, A2 => n4791, B1 => N12285, B2 => 
                           n305, ZN => n4824);
   U5431 : OAI21_X1 port map( B1 => n11830, B2 => n4789, A => n4825, ZN => 
                           n13173);
   U5432 : AOI22_X1 port map( A1 => N13848, A2 => n4791, B1 => N12286, B2 => 
                           n305, ZN => n4825);
   U5433 : OAI21_X1 port map( B1 => n11829, B2 => n4789, A => n4826, ZN => 
                           n13172);
   U5434 : AOI22_X1 port map( A1 => N13849, A2 => n4791, B1 => N12287, B2 => 
                           n305, ZN => n4826);
   U5435 : OAI21_X1 port map( B1 => n11828, B2 => n4789, A => n4827, ZN => 
                           n13171);
   U5436 : AOI22_X1 port map( A1 => N13850, A2 => n4791, B1 => N12288, B2 => 
                           n305, ZN => n4827);
   U5437 : OAI21_X1 port map( B1 => n11827, B2 => n4789, A => n4828, ZN => 
                           n13170);
   U5438 : AOI22_X1 port map( A1 => N13851, A2 => n4791, B1 => N12289, B2 => 
                           n305, ZN => n4828);
   U5439 : OAI21_X1 port map( B1 => n11826, B2 => n4789, A => n4829, ZN => 
                           n13169);
   U5440 : AOI22_X1 port map( A1 => N13852, A2 => n4791, B1 => N12290, B2 => 
                           n305, ZN => n4829);
   U5441 : OAI21_X1 port map( B1 => n11825, B2 => n4789, A => n4830, ZN => 
                           n13168);
   U5442 : AOI22_X1 port map( A1 => N13853, A2 => n4791, B1 => N12291, B2 => 
                           n305, ZN => n4830);
   U5443 : OAI21_X1 port map( B1 => n11824, B2 => n4789, A => n4831, ZN => 
                           n13167);
   U5444 : AOI22_X1 port map( A1 => N13854, A2 => n4791, B1 => N12292, B2 => 
                           n305, ZN => n4831);
   U5445 : OAI21_X1 port map( B1 => n11823, B2 => n4789, A => n4832, ZN => 
                           n13166);
   U5446 : AOI22_X1 port map( A1 => N13855, A2 => n4791, B1 => N12293, B2 => 
                           n305, ZN => n4832);
   U5447 : OAI21_X1 port map( B1 => n11822, B2 => n4789, A => n4833, ZN => 
                           n13165);
   U5448 : AOI22_X1 port map( A1 => N13856, A2 => n4791, B1 => N12294, B2 => 
                           n305, ZN => n4833);
   U5449 : OAI21_X1 port map( B1 => n11821, B2 => n4789, A => n4834, ZN => 
                           n13164);
   U5450 : AOI22_X1 port map( A1 => N13857, A2 => n4791, B1 => N12295, B2 => 
                           n305, ZN => n4834);
   U5451 : OAI21_X1 port map( B1 => n11820, B2 => n4789, A => n4835, ZN => 
                           n13163);
   U5452 : AOI22_X1 port map( A1 => N13858, A2 => n4791, B1 => N12296, B2 => 
                           n305, ZN => n4835);
   U5453 : OAI21_X1 port map( B1 => n11819, B2 => n4789, A => n4836, ZN => 
                           n13162);
   U5454 : AOI22_X1 port map( A1 => N13859, A2 => n4791, B1 => N12297, B2 => 
                           n305, ZN => n4836);
   U5455 : OAI21_X1 port map( B1 => n11818, B2 => n4789, A => n4837, ZN => 
                           n13161);
   U5456 : AOI22_X1 port map( A1 => N13860, A2 => n4791, B1 => N12298, B2 => 
                           n305, ZN => n4837);
   U5457 : OAI21_X1 port map( B1 => n11817, B2 => n4789, A => n4838, ZN => 
                           n13160);
   U5458 : AOI22_X1 port map( A1 => N13861, A2 => n4791, B1 => N12299, B2 => 
                           n305, ZN => n4838);
   U5459 : AOI22_X1 port map( A1 => CALL, A2 => n16455, B1 => n4840, B2 => 
                           n4784, ZN => n4802);
   U5460 : INV_X1 port map( A => n4811, ZN => n4808);
   U5461 : NAND2_X1 port map( A1 => n4789, A2 => n4841, ZN => n4839);
   U5462 : NAND2_X1 port map( A1 => ENABLE, A2 => n4842, ZN => n4800);
   U5463 : NAND3_X1 port map( A1 => n4843, A2 => n4844, A3 => n4845, ZN => 
                           n4842);
   U5464 : NOR3_X1 port map( A1 => n4811, A2 => RESET, A3 => n4812, ZN => n4845
                           );
   U5465 : NOR3_X1 port map( A1 => n4846, A2 => n16455, A3 => n4847, ZN => 
                           n4811);
   U5466 : NAND2_X1 port map( A1 => n4848, A2 => n4849, ZN => n13159);
   U5467 : NAND3_X1 port map( A1 => CALL, A2 => n4850, A3 => ENABLE, ZN => 
                           n4849);
   U5468 : OAI21_X1 port map( B1 => n4786, B2 => n4850, A => n117, ZN => n4848)
                           ;
   U5469 : NAND3_X1 port map( A1 => RET, A2 => n116, A3 => n4810, ZN => n4850);
   U5470 : OAI21_X1 port map( B1 => n11869, B2 => n210, A => n4852, ZN => 
                           n13158);
   U5471 : AOI22_X1 port map( A1 => N50337, A2 => n207, B1 => N12237, B2 => 
                           n214, ZN => n4852);
   U5472 : OAI21_X1 port map( B1 => n11868, B2 => n210, A => n4853, ZN => 
                           n13157);
   U5473 : AOI22_X1 port map( A1 => N50338, A2 => n207, B1 => N12238, B2 => 
                           n214, ZN => n4853);
   U5474 : NAND2_X1 port map( A1 => n4854, A2 => n4855, ZN => n13156);
   U5475 : OAI211_X1 port map( C1 => n4784, C2 => N12239, A => n210, B => n4809
                           , ZN => n4855);
   U5476 : OAI21_X1 port map( B1 => n207, B2 => n209, A => n1, ZN => n4854);
   U5477 : OAI21_X1 port map( B1 => n11866, B2 => n210, A => n4856, ZN => 
                           n13155);
   U5478 : AOI22_X1 port map( A1 => N50340, A2 => n207, B1 => N12240, B2 => 
                           n214, ZN => n4856);
   U5479 : OAI21_X1 port map( B1 => n11865, B2 => n210, A => n4857, ZN => 
                           n13154);
   U5480 : AOI22_X1 port map( A1 => N50341, A2 => n207, B1 => N12241, B2 => 
                           n214, ZN => n4857);
   U5481 : OAI21_X1 port map( B1 => n11864, B2 => n210, A => n4858, ZN => 
                           n13153);
   U5482 : AOI22_X1 port map( A1 => N50342, A2 => n207, B1 => N12242, B2 => 
                           n214, ZN => n4858);
   U5483 : NAND3_X1 port map( A1 => n4859, A2 => n4860, A3 => n4861, ZN => 
                           n13152);
   U5484 : AOI221_X1 port map( B1 => n4862, B2 => n4863, C1 => MEM_IN(0), C2 =>
                           n206, A => n4864, ZN => n4861);
   U5485 : OAI22_X1 port map( A1 => n11789, A2 => n4865, B1 => n4866, B2 => 
                           n4867, ZN => n4864);
   U5486 : AOI22_X1 port map( A1 => n4868, A2 => n4869, B1 => n4870, B2 => 
                           n4871, ZN => n4860);
   U5487 : AOI22_X1 port map( A1 => n4872, A2 => n4873, B1 => n4874, B2 => 
                           n4875, ZN => n4859);
   U5488 : NAND3_X1 port map( A1 => n4876, A2 => n4877, A3 => n4878, ZN => 
                           n13151);
   U5489 : AOI221_X1 port map( B1 => n4879, B2 => n4862, C1 => MEM_IN(1), C2 =>
                           n206, A => n4880, ZN => n4878);
   U5490 : OAI22_X1 port map( A1 => n11788, A2 => n4865, B1 => n4866, B2 => 
                           n4881, ZN => n4880);
   U5491 : AOI22_X1 port map( A1 => n4868, A2 => n4882, B1 => n4870, B2 => 
                           n4883, ZN => n4877);
   U5492 : AOI22_X1 port map( A1 => n4872, A2 => n4884, B1 => n4874, B2 => 
                           n4885, ZN => n4876);
   U5493 : NAND3_X1 port map( A1 => n4886, A2 => n4887, A3 => n4888, ZN => 
                           n13150);
   U5494 : AOI221_X1 port map( B1 => n4889, B2 => n4862, C1 => MEM_IN(2), C2 =>
                           n206, A => n4890, ZN => n4888);
   U5495 : OAI22_X1 port map( A1 => n11787, A2 => n4865, B1 => n4866, B2 => 
                           n4891, ZN => n4890);
   U5496 : AOI22_X1 port map( A1 => n4868, A2 => n4892, B1 => n4870, B2 => 
                           n4893, ZN => n4887);
   U5497 : AOI22_X1 port map( A1 => n4872, A2 => n4894, B1 => n4874, B2 => 
                           n4895, ZN => n4886);
   U5498 : NAND3_X1 port map( A1 => n4896, A2 => n4897, A3 => n4898, ZN => 
                           n13149);
   U5499 : AOI221_X1 port map( B1 => n4899, B2 => n4862, C1 => MEM_IN(3), C2 =>
                           n206, A => n4900, ZN => n4898);
   U5500 : OAI22_X1 port map( A1 => n11786, A2 => n4865, B1 => n4866, B2 => 
                           n4901, ZN => n4900);
   U5501 : AOI22_X1 port map( A1 => n4868, A2 => n4902, B1 => n4870, B2 => 
                           n4903, ZN => n4897);
   U5502 : AOI22_X1 port map( A1 => n4872, A2 => n4904, B1 => n4874, B2 => 
                           n4905, ZN => n4896);
   U5503 : NAND3_X1 port map( A1 => n4906, A2 => n4907, A3 => n4908, ZN => 
                           n13148);
   U5504 : AOI221_X1 port map( B1 => n4909, B2 => n4862, C1 => MEM_IN(4), C2 =>
                           n206, A => n4910, ZN => n4908);
   U5505 : OAI22_X1 port map( A1 => n11785, A2 => n4865, B1 => n4866, B2 => 
                           n4911, ZN => n4910);
   U5506 : AOI22_X1 port map( A1 => n4868, A2 => n4912, B1 => n4870, B2 => 
                           n4913, ZN => n4907);
   U5507 : AOI22_X1 port map( A1 => n4872, A2 => n4914, B1 => n4874, B2 => 
                           n4915, ZN => n4906);
   U5508 : NAND3_X1 port map( A1 => n4916, A2 => n4917, A3 => n4918, ZN => 
                           n13147);
   U5509 : AOI221_X1 port map( B1 => n4919, B2 => n4862, C1 => MEM_IN(5), C2 =>
                           n206, A => n4920, ZN => n4918);
   U5510 : OAI22_X1 port map( A1 => n11784, A2 => n4865, B1 => n4866, B2 => 
                           n4921, ZN => n4920);
   U5511 : AOI22_X1 port map( A1 => n4868, A2 => n4922, B1 => n4870, B2 => 
                           n4923, ZN => n4917);
   U5512 : AOI22_X1 port map( A1 => n4872, A2 => n4924, B1 => n4874, B2 => 
                           n4925, ZN => n4916);
   U5513 : NAND3_X1 port map( A1 => n4926, A2 => n4927, A3 => n4928, ZN => 
                           n13146);
   U5514 : AOI221_X1 port map( B1 => n4929, B2 => n4862, C1 => MEM_IN(6), C2 =>
                           n206, A => n4930, ZN => n4928);
   U5515 : OAI22_X1 port map( A1 => n11783, A2 => n4865, B1 => n4866, B2 => 
                           n4931, ZN => n4930);
   U5516 : AOI22_X1 port map( A1 => n4868, A2 => n4932, B1 => n4870, B2 => 
                           n4933, ZN => n4927);
   U5517 : AOI22_X1 port map( A1 => n4872, A2 => n4934, B1 => n4874, B2 => 
                           n4935, ZN => n4926);
   U5518 : NAND3_X1 port map( A1 => n4936, A2 => n4937, A3 => n4938, ZN => 
                           n13145);
   U5519 : AOI221_X1 port map( B1 => n4939, B2 => n4862, C1 => MEM_IN(7), C2 =>
                           n206, A => n4940, ZN => n4938);
   U5520 : OAI22_X1 port map( A1 => n11782, A2 => n4865, B1 => n4866, B2 => 
                           n4941, ZN => n4940);
   U5521 : AOI22_X1 port map( A1 => n4868, A2 => n4942, B1 => n4870, B2 => 
                           n4943, ZN => n4937);
   U5522 : AOI22_X1 port map( A1 => n4872, A2 => n4944, B1 => n4874, B2 => 
                           n4945, ZN => n4936);
   U5523 : NAND3_X1 port map( A1 => n4946, A2 => n4947, A3 => n4948, ZN => 
                           n13144);
   U5524 : AOI221_X1 port map( B1 => n4949, B2 => n4862, C1 => MEM_IN(8), C2 =>
                           n206, A => n4950, ZN => n4948);
   U5525 : OAI22_X1 port map( A1 => n11781, A2 => n4865, B1 => n4866, B2 => 
                           n4951, ZN => n4950);
   U5526 : AOI22_X1 port map( A1 => n4868, A2 => n4952, B1 => n4870, B2 => 
                           n4953, ZN => n4947);
   U5527 : AOI22_X1 port map( A1 => n4872, A2 => n4954, B1 => n4874, B2 => 
                           n4955, ZN => n4946);
   U5528 : NAND3_X1 port map( A1 => n4956, A2 => n4957, A3 => n4958, ZN => 
                           n13143);
   U5529 : AOI221_X1 port map( B1 => n4959, B2 => n4862, C1 => MEM_IN(9), C2 =>
                           n206, A => n4960, ZN => n4958);
   U5530 : OAI22_X1 port map( A1 => n11780, A2 => n4865, B1 => n4866, B2 => 
                           n4961, ZN => n4960);
   U5531 : AOI22_X1 port map( A1 => n4868, A2 => n4962, B1 => n4870, B2 => 
                           n4963, ZN => n4957);
   U5532 : AOI22_X1 port map( A1 => n4872, A2 => n4964, B1 => n4874, B2 => 
                           n4965, ZN => n4956);
   U5533 : NAND3_X1 port map( A1 => n4966, A2 => n4967, A3 => n4968, ZN => 
                           n13142);
   U5534 : AOI221_X1 port map( B1 => n4969, B2 => n4862, C1 => MEM_IN(10), C2 
                           => n206, A => n4970, ZN => n4968);
   U5535 : OAI22_X1 port map( A1 => n11779, A2 => n4865, B1 => n4866, B2 => 
                           n4971, ZN => n4970);
   U5536 : AOI22_X1 port map( A1 => n4868, A2 => n4972, B1 => n4870, B2 => 
                           n4973, ZN => n4967);
   U5537 : AOI22_X1 port map( A1 => n4872, A2 => n4974, B1 => n4874, B2 => 
                           n4975, ZN => n4966);
   U5538 : NAND3_X1 port map( A1 => n4976, A2 => n4977, A3 => n4978, ZN => 
                           n13141);
   U5539 : AOI221_X1 port map( B1 => n4979, B2 => n4862, C1 => MEM_IN(11), C2 
                           => n206, A => n4980, ZN => n4978);
   U5540 : OAI22_X1 port map( A1 => n11778, A2 => n4865, B1 => n4866, B2 => 
                           n4981, ZN => n4980);
   U5541 : AOI22_X1 port map( A1 => n4868, A2 => n4982, B1 => n4870, B2 => 
                           n4983, ZN => n4977);
   U5542 : AOI22_X1 port map( A1 => n4872, A2 => n4984, B1 => n4874, B2 => 
                           n4985, ZN => n4976);
   U5543 : NAND3_X1 port map( A1 => n4986, A2 => n4987, A3 => n4988, ZN => 
                           n13140);
   U5544 : AOI221_X1 port map( B1 => n4989, B2 => n4862, C1 => MEM_IN(12), C2 
                           => n206, A => n4990, ZN => n4988);
   U5545 : OAI22_X1 port map( A1 => n11777, A2 => n4865, B1 => n4866, B2 => 
                           n4991, ZN => n4990);
   U5546 : AOI22_X1 port map( A1 => n4868, A2 => n4992, B1 => n4870, B2 => 
                           n4993, ZN => n4987);
   U5547 : AOI22_X1 port map( A1 => n4872, A2 => n4994, B1 => n4874, B2 => 
                           n4995, ZN => n4986);
   U5548 : NAND3_X1 port map( A1 => n4996, A2 => n4997, A3 => n4998, ZN => 
                           n13139);
   U5549 : AOI221_X1 port map( B1 => n4999, B2 => n4862, C1 => MEM_IN(13), C2 
                           => n206, A => n5000, ZN => n4998);
   U5550 : OAI22_X1 port map( A1 => n11776, A2 => n4865, B1 => n4866, B2 => 
                           n5001, ZN => n5000);
   U5551 : AOI22_X1 port map( A1 => n4868, A2 => n5002, B1 => n4870, B2 => 
                           n5003, ZN => n4997);
   U5552 : AOI22_X1 port map( A1 => n4872, A2 => n5004, B1 => n4874, B2 => 
                           n5005, ZN => n4996);
   U5553 : NAND3_X1 port map( A1 => n5006, A2 => n5007, A3 => n5008, ZN => 
                           n13138);
   U5554 : AOI221_X1 port map( B1 => n5009, B2 => n4862, C1 => MEM_IN(14), C2 
                           => n206, A => n5010, ZN => n5008);
   U5555 : OAI22_X1 port map( A1 => n11775, A2 => n4865, B1 => n4866, B2 => 
                           n5011, ZN => n5010);
   U5556 : AOI22_X1 port map( A1 => n4868, A2 => n5012, B1 => n4870, B2 => 
                           n5013, ZN => n5007);
   U5557 : AOI22_X1 port map( A1 => n4872, A2 => n5014, B1 => n4874, B2 => 
                           n5015, ZN => n5006);
   U5558 : NAND3_X1 port map( A1 => n5016, A2 => n5017, A3 => n5018, ZN => 
                           n13137);
   U5559 : AOI221_X1 port map( B1 => n5019, B2 => n4862, C1 => MEM_IN(15), C2 
                           => n206, A => n5020, ZN => n5018);
   U5560 : OAI22_X1 port map( A1 => n11774, A2 => n4865, B1 => n4866, B2 => 
                           n5021, ZN => n5020);
   U5561 : AOI22_X1 port map( A1 => n4868, A2 => n5022, B1 => n4870, B2 => 
                           n5023, ZN => n5017);
   U5562 : AOI22_X1 port map( A1 => n4872, A2 => n5024, B1 => n4874, B2 => 
                           n5025, ZN => n5016);
   U5563 : NAND3_X1 port map( A1 => n5026, A2 => n5027, A3 => n5028, ZN => 
                           n13136);
   U5564 : AOI221_X1 port map( B1 => n5029, B2 => n4862, C1 => MEM_IN(16), C2 
                           => n206, A => n5030, ZN => n5028);
   U5565 : OAI22_X1 port map( A1 => n11773, A2 => n4865, B1 => n4866, B2 => 
                           n5031, ZN => n5030);
   U5566 : AOI22_X1 port map( A1 => n4868, A2 => n5032, B1 => n4870, B2 => 
                           n5033, ZN => n5027);
   U5567 : AOI22_X1 port map( A1 => n4872, A2 => n5034, B1 => n4874, B2 => 
                           n5035, ZN => n5026);
   U5568 : NAND3_X1 port map( A1 => n5036, A2 => n5037, A3 => n5038, ZN => 
                           n13135);
   U5569 : AOI221_X1 port map( B1 => n5039, B2 => n4862, C1 => MEM_IN(17), C2 
                           => n206, A => n5040, ZN => n5038);
   U5570 : OAI22_X1 port map( A1 => n11772, A2 => n4865, B1 => n4866, B2 => 
                           n5041, ZN => n5040);
   U5571 : AOI22_X1 port map( A1 => n4868, A2 => n5042, B1 => n4870, B2 => 
                           n5043, ZN => n5037);
   U5572 : AOI22_X1 port map( A1 => n4872, A2 => n5044, B1 => n4874, B2 => 
                           n5045, ZN => n5036);
   U5573 : NAND3_X1 port map( A1 => n5046, A2 => n5047, A3 => n5048, ZN => 
                           n13134);
   U5574 : AOI221_X1 port map( B1 => n5049, B2 => n4862, C1 => MEM_IN(18), C2 
                           => n206, A => n5050, ZN => n5048);
   U5575 : OAI22_X1 port map( A1 => n11771, A2 => n4865, B1 => n4866, B2 => 
                           n5051, ZN => n5050);
   U5576 : AOI22_X1 port map( A1 => n4868, A2 => n5052, B1 => n4870, B2 => 
                           n5053, ZN => n5047);
   U5577 : AOI22_X1 port map( A1 => n4872, A2 => n5054, B1 => n4874, B2 => 
                           n5055, ZN => n5046);
   U5578 : NAND3_X1 port map( A1 => n5056, A2 => n5057, A3 => n5058, ZN => 
                           n13133);
   U5579 : AOI221_X1 port map( B1 => n5059, B2 => n4862, C1 => MEM_IN(19), C2 
                           => n206, A => n5060, ZN => n5058);
   U5580 : OAI22_X1 port map( A1 => n11770, A2 => n4865, B1 => n4866, B2 => 
                           n5061, ZN => n5060);
   U5581 : AOI22_X1 port map( A1 => n4868, A2 => n5062, B1 => n4870, B2 => 
                           n5063, ZN => n5057);
   U5582 : AOI22_X1 port map( A1 => n4872, A2 => n5064, B1 => n4874, B2 => 
                           n5065, ZN => n5056);
   U5583 : NAND3_X1 port map( A1 => n5066, A2 => n5067, A3 => n5068, ZN => 
                           n13132);
   U5584 : AOI221_X1 port map( B1 => n5069, B2 => n4862, C1 => MEM_IN(20), C2 
                           => n206, A => n5070, ZN => n5068);
   U5585 : OAI22_X1 port map( A1 => n11769, A2 => n4865, B1 => n4866, B2 => 
                           n5071, ZN => n5070);
   U5586 : AOI22_X1 port map( A1 => n4868, A2 => n5072, B1 => n4870, B2 => 
                           n5073, ZN => n5067);
   U5587 : AOI22_X1 port map( A1 => n4872, A2 => n5074, B1 => n4874, B2 => 
                           n5075, ZN => n5066);
   U5588 : NAND3_X1 port map( A1 => n5076, A2 => n5077, A3 => n5078, ZN => 
                           n13131);
   U5589 : AOI221_X1 port map( B1 => n5079, B2 => n4862, C1 => MEM_IN(21), C2 
                           => n206, A => n5080, ZN => n5078);
   U5590 : OAI22_X1 port map( A1 => n11768, A2 => n4865, B1 => n4866, B2 => 
                           n5081, ZN => n5080);
   U5591 : AOI22_X1 port map( A1 => n4868, A2 => n5082, B1 => n4870, B2 => 
                           n5083, ZN => n5077);
   U5592 : AOI22_X1 port map( A1 => n4872, A2 => n5084, B1 => n4874, B2 => 
                           n5085, ZN => n5076);
   U5593 : NAND3_X1 port map( A1 => n5086, A2 => n5087, A3 => n5088, ZN => 
                           n13130);
   U5594 : AOI221_X1 port map( B1 => n5089, B2 => n4862, C1 => MEM_IN(22), C2 
                           => n206, A => n5090, ZN => n5088);
   U5595 : OAI22_X1 port map( A1 => n11767, A2 => n4865, B1 => n4866, B2 => 
                           n5091, ZN => n5090);
   U5596 : AOI22_X1 port map( A1 => n4868, A2 => n5092, B1 => n4870, B2 => 
                           n5093, ZN => n5087);
   U5597 : AOI22_X1 port map( A1 => n4872, A2 => n5094, B1 => n4874, B2 => 
                           n5095, ZN => n5086);
   U5598 : NAND3_X1 port map( A1 => n5096, A2 => n5097, A3 => n5098, ZN => 
                           n13129);
   U5599 : AOI221_X1 port map( B1 => n5099, B2 => n4862, C1 => MEM_IN(23), C2 
                           => n206, A => n5100, ZN => n5098);
   U5600 : OAI22_X1 port map( A1 => n11766, A2 => n4865, B1 => n4866, B2 => 
                           n5101, ZN => n5100);
   U5601 : AOI22_X1 port map( A1 => n4868, A2 => n5102, B1 => n4870, B2 => 
                           n5103, ZN => n5097);
   U5602 : AOI22_X1 port map( A1 => n4872, A2 => n5104, B1 => n4874, B2 => 
                           n5105, ZN => n5096);
   U5603 : NAND3_X1 port map( A1 => n5106, A2 => n5107, A3 => n5108, ZN => 
                           n13128);
   U5604 : AOI221_X1 port map( B1 => n5109, B2 => n4862, C1 => MEM_IN(24), C2 
                           => n206, A => n5110, ZN => n5108);
   U5605 : OAI22_X1 port map( A1 => n11765, A2 => n4865, B1 => n4866, B2 => 
                           n5111, ZN => n5110);
   U5606 : AOI22_X1 port map( A1 => n4868, A2 => n5112, B1 => n4870, B2 => 
                           n5113, ZN => n5107);
   U5607 : AOI22_X1 port map( A1 => n4872, A2 => n5114, B1 => n4874, B2 => 
                           n5115, ZN => n5106);
   U5608 : NAND3_X1 port map( A1 => n5116, A2 => n5117, A3 => n5118, ZN => 
                           n13127);
   U5609 : AOI221_X1 port map( B1 => n5119, B2 => n4862, C1 => MEM_IN(25), C2 
                           => n206, A => n5120, ZN => n5118);
   U5610 : OAI22_X1 port map( A1 => n11764, A2 => n4865, B1 => n4866, B2 => 
                           n5121, ZN => n5120);
   U5611 : AOI22_X1 port map( A1 => n4868, A2 => n5122, B1 => n4870, B2 => 
                           n5123, ZN => n5117);
   U5612 : AOI22_X1 port map( A1 => n4872, A2 => n5124, B1 => n4874, B2 => 
                           n5125, ZN => n5116);
   U5613 : NAND3_X1 port map( A1 => n5126, A2 => n5127, A3 => n5128, ZN => 
                           n13126);
   U5614 : AOI221_X1 port map( B1 => n5129, B2 => n4862, C1 => MEM_IN(26), C2 
                           => n206, A => n5130, ZN => n5128);
   U5615 : OAI22_X1 port map( A1 => n11763, A2 => n4865, B1 => n4866, B2 => 
                           n5131, ZN => n5130);
   U5616 : AOI22_X1 port map( A1 => n4868, A2 => n5132, B1 => n4870, B2 => 
                           n5133, ZN => n5127);
   U5617 : AOI22_X1 port map( A1 => n4872, A2 => n5134, B1 => n4874, B2 => 
                           n5135, ZN => n5126);
   U5618 : NAND3_X1 port map( A1 => n5136, A2 => n5137, A3 => n5138, ZN => 
                           n13125);
   U5619 : AOI221_X1 port map( B1 => n5139, B2 => n4862, C1 => MEM_IN(27), C2 
                           => n206, A => n5140, ZN => n5138);
   U5620 : OAI22_X1 port map( A1 => n11762, A2 => n4865, B1 => n4866, B2 => 
                           n5141, ZN => n5140);
   U5621 : AOI22_X1 port map( A1 => n4868, A2 => n5142, B1 => n4870, B2 => 
                           n5143, ZN => n5137);
   U5622 : AOI22_X1 port map( A1 => n4872, A2 => n5144, B1 => n4874, B2 => 
                           n5145, ZN => n5136);
   U5623 : NAND3_X1 port map( A1 => n5146, A2 => n5147, A3 => n5148, ZN => 
                           n13124);
   U5624 : AOI221_X1 port map( B1 => n5149, B2 => n4862, C1 => MEM_IN(28), C2 
                           => n206, A => n5150, ZN => n5148);
   U5625 : OAI22_X1 port map( A1 => n11761, A2 => n4865, B1 => n4866, B2 => 
                           n5151, ZN => n5150);
   U5626 : AOI22_X1 port map( A1 => n4868, A2 => n5152, B1 => n4870, B2 => 
                           n5153, ZN => n5147);
   U5627 : AOI22_X1 port map( A1 => n4872, A2 => n5154, B1 => n4874, B2 => 
                           n5155, ZN => n5146);
   U5628 : NAND3_X1 port map( A1 => n5156, A2 => n5157, A3 => n5158, ZN => 
                           n13123);
   U5629 : AOI221_X1 port map( B1 => n5159, B2 => n4862, C1 => MEM_IN(29), C2 
                           => n206, A => n5160, ZN => n5158);
   U5630 : OAI22_X1 port map( A1 => n11760, A2 => n4865, B1 => n4866, B2 => 
                           n5161, ZN => n5160);
   U5631 : AOI22_X1 port map( A1 => n4868, A2 => n5162, B1 => n4870, B2 => 
                           n5163, ZN => n5157);
   U5632 : AOI22_X1 port map( A1 => n4872, A2 => n5164, B1 => n4874, B2 => 
                           n5165, ZN => n5156);
   U5633 : NAND3_X1 port map( A1 => n5166, A2 => n5167, A3 => n5168, ZN => 
                           n13122);
   U5634 : AOI221_X1 port map( B1 => n5169, B2 => n4862, C1 => MEM_IN(30), C2 
                           => n206, A => n5170, ZN => n5168);
   U5635 : OAI22_X1 port map( A1 => n11759, A2 => n4865, B1 => n4866, B2 => 
                           n5171, ZN => n5170);
   U5636 : AOI22_X1 port map( A1 => n4868, A2 => n5172, B1 => n4870, B2 => 
                           n5173, ZN => n5167);
   U5637 : AOI22_X1 port map( A1 => n4872, A2 => n5174, B1 => n4874, B2 => 
                           n5175, ZN => n5166);
   U5638 : NAND3_X1 port map( A1 => n5176, A2 => n5177, A3 => n5178, ZN => 
                           n13121);
   U5639 : AOI221_X1 port map( B1 => n5179, B2 => n4862, C1 => MEM_IN(31), C2 
                           => n206, A => n5180, ZN => n5178);
   U5640 : OAI22_X1 port map( A1 => n11758, A2 => n4865, B1 => n4866, B2 => 
                           n5181, ZN => n5180);
   U5641 : OAI21_X1 port map( B1 => n5186, B2 => n4787, A => n5187, ZN => n5185
                           );
   U5642 : NOR3_X1 port map( A1 => n5188, A2 => n5189, A3 => n5190, ZN => n5186
                           );
   U5643 : AOI22_X1 port map( A1 => n4868, A2 => n5191, B1 => n4870, B2 => 
                           n5192, ZN => n5177);
   U5644 : AOI22_X1 port map( A1 => n4872, A2 => n5195, B1 => n4874, B2 => 
                           n5196, ZN => n5176);
   U5645 : OAI22_X1 port map( A1 => n5199, A2 => n5183, B1 => n208, B2 => n5200
                           , ZN => n5187);
   U5646 : INV_X1 port map( A => n4865, ZN => n5200);
   U5647 : NAND3_X1 port map( A1 => n5201, A2 => n4865, A3 => n208, ZN => n5183
                           );
   U5648 : NAND3_X1 port map( A1 => n5206, A2 => ENABLE, A3 => n5189, ZN => 
                           n5205);
   U5649 : NOR2_X1 port map( A1 => n5182, A2 => n5199, ZN => n5203);
   U5650 : INV_X1 port map( A => n5201, ZN => n5182);
   U5651 : AOI21_X1 port map( B1 => n5207, B2 => n5208, A => n5209, ZN => n5202
                           );
   U5652 : NOR3_X1 port map( A1 => n5210, A2 => n5189, A3 => n5211, ZN => n5201
                           );
   U5653 : INV_X1 port map( A => n5212, ZN => n5210);
   U5654 : INV_X1 port map( A => n5184, ZN => n5199);
   U5655 : NOR2_X1 port map( A1 => n5213, A2 => n5214, ZN => n5184);
   U5656 : AND2_X1 port map( A1 => n5215, A2 => n5216, ZN => n5189);
   U5657 : NAND3_X1 port map( A1 => n5217, A2 => n5218, A3 => n5219, ZN => 
                           n13120);
   U5658 : AOI221_X1 port map( B1 => n5220, B2 => n4863, C1 => n5221, C2 => 
                           MEM_IN(0), A => n5222, ZN => n5219);
   U5659 : OAI22_X1 port map( A1 => n11757, A2 => n231, B1 => n4867, B2 => 
                           n5224, ZN => n5222);
   U5660 : AOI22_X1 port map( A1 => n5225, A2 => n4869, B1 => n5226, B2 => 
                           n4871, ZN => n5218);
   U5661 : AOI22_X1 port map( A1 => n5227, A2 => n4873, B1 => n5228, B2 => 
                           n4875, ZN => n5217);
   U5662 : NAND3_X1 port map( A1 => n5229, A2 => n5230, A3 => n5231, ZN => 
                           n13119);
   U5663 : AOI221_X1 port map( B1 => n5220, B2 => n4879, C1 => n5221, C2 => 
                           MEM_IN(1), A => n5232, ZN => n5231);
   U5664 : OAI22_X1 port map( A1 => n11756, A2 => n231, B1 => n4881, B2 => 
                           n5224, ZN => n5232);
   U5665 : AOI22_X1 port map( A1 => n5225, A2 => n4882, B1 => n5226, B2 => 
                           n4883, ZN => n5230);
   U5666 : AOI22_X1 port map( A1 => n5227, A2 => n4884, B1 => n5228, B2 => 
                           n4885, ZN => n5229);
   U5667 : NAND3_X1 port map( A1 => n5233, A2 => n5234, A3 => n5235, ZN => 
                           n13118);
   U5668 : AOI221_X1 port map( B1 => n5220, B2 => n4889, C1 => n5221, C2 => 
                           MEM_IN(2), A => n5236, ZN => n5235);
   U5669 : OAI22_X1 port map( A1 => n11755, A2 => n231, B1 => n4891, B2 => 
                           n5224, ZN => n5236);
   U5670 : AOI22_X1 port map( A1 => n5225, A2 => n4892, B1 => n5226, B2 => 
                           n4893, ZN => n5234);
   U5671 : AOI22_X1 port map( A1 => n5227, A2 => n4894, B1 => n5228, B2 => 
                           n4895, ZN => n5233);
   U5672 : NAND3_X1 port map( A1 => n5237, A2 => n5238, A3 => n5239, ZN => 
                           n13117);
   U5673 : AOI221_X1 port map( B1 => n5220, B2 => n4899, C1 => n5221, C2 => 
                           MEM_IN(3), A => n5240, ZN => n5239);
   U5674 : OAI22_X1 port map( A1 => n11754, A2 => n231, B1 => n4901, B2 => 
                           n5224, ZN => n5240);
   U5675 : AOI22_X1 port map( A1 => n5225, A2 => n4902, B1 => n5226, B2 => 
                           n4903, ZN => n5238);
   U5676 : AOI22_X1 port map( A1 => n5227, A2 => n4904, B1 => n5228, B2 => 
                           n4905, ZN => n5237);
   U5677 : NAND3_X1 port map( A1 => n5241, A2 => n5242, A3 => n5243, ZN => 
                           n13116);
   U5678 : AOI221_X1 port map( B1 => n5220, B2 => n4909, C1 => n5221, C2 => 
                           MEM_IN(4), A => n5244, ZN => n5243);
   U5679 : OAI22_X1 port map( A1 => n11753, A2 => n231, B1 => n4911, B2 => 
                           n5224, ZN => n5244);
   U5680 : AOI22_X1 port map( A1 => n5225, A2 => n4912, B1 => n5226, B2 => 
                           n4913, ZN => n5242);
   U5681 : AOI22_X1 port map( A1 => n5227, A2 => n4914, B1 => n5228, B2 => 
                           n4915, ZN => n5241);
   U5682 : NAND3_X1 port map( A1 => n5245, A2 => n5246, A3 => n5247, ZN => 
                           n13115);
   U5683 : AOI221_X1 port map( B1 => n5220, B2 => n4919, C1 => n5221, C2 => 
                           MEM_IN(5), A => n5248, ZN => n5247);
   U5684 : OAI22_X1 port map( A1 => n11752, A2 => n231, B1 => n4921, B2 => 
                           n5224, ZN => n5248);
   U5685 : AOI22_X1 port map( A1 => n5225, A2 => n4922, B1 => n5226, B2 => 
                           n4923, ZN => n5246);
   U5686 : AOI22_X1 port map( A1 => n5227, A2 => n4924, B1 => n5228, B2 => 
                           n4925, ZN => n5245);
   U5687 : NAND3_X1 port map( A1 => n5249, A2 => n5250_port, A3 => n5251_port, 
                           ZN => n13114);
   U5688 : AOI221_X1 port map( B1 => n5220, B2 => n4929, C1 => n5221, C2 => 
                           MEM_IN(6), A => n5252_port, ZN => n5251_port);
   U5689 : OAI22_X1 port map( A1 => n11751, A2 => n231, B1 => n4931, B2 => 
                           n5224, ZN => n5252_port);
   U5690 : AOI22_X1 port map( A1 => n5225, A2 => n4932, B1 => n5226, B2 => 
                           n4933, ZN => n5250_port);
   U5691 : AOI22_X1 port map( A1 => n5227, A2 => n4934, B1 => n5228, B2 => 
                           n4935, ZN => n5249);
   U5692 : NAND3_X1 port map( A1 => n5253_port, A2 => n5254_port, A3 => 
                           n5255_port, ZN => n13113);
   U5693 : AOI221_X1 port map( B1 => n5220, B2 => n4939, C1 => n5221, C2 => 
                           MEM_IN(7), A => n5256_port, ZN => n5255_port);
   U5694 : OAI22_X1 port map( A1 => n11750, A2 => n231, B1 => n4941, B2 => 
                           n5224, ZN => n5256_port);
   U5695 : AOI22_X1 port map( A1 => n5225, A2 => n4942, B1 => n5226, B2 => 
                           n4943, ZN => n5254_port);
   U5696 : AOI22_X1 port map( A1 => n5227, A2 => n4944, B1 => n5228, B2 => 
                           n4945, ZN => n5253_port);
   U5697 : NAND3_X1 port map( A1 => n5257_port, A2 => n5258_port, A3 => 
                           n5259_port, ZN => n13112);
   U5698 : AOI221_X1 port map( B1 => n5220, B2 => n4949, C1 => n5221, C2 => 
                           MEM_IN(8), A => n5260_port, ZN => n5259_port);
   U5699 : OAI22_X1 port map( A1 => n11749, A2 => n231, B1 => n4951, B2 => 
                           n5224, ZN => n5260_port);
   U5700 : AOI22_X1 port map( A1 => n5225, A2 => n4952, B1 => n5226, B2 => 
                           n4953, ZN => n5258_port);
   U5701 : AOI22_X1 port map( A1 => n5227, A2 => n4954, B1 => n5228, B2 => 
                           n4955, ZN => n5257_port);
   U5702 : NAND3_X1 port map( A1 => n5261_port, A2 => n5262_port, A3 => 
                           n5263_port, ZN => n13111);
   U5703 : AOI221_X1 port map( B1 => n5220, B2 => n4959, C1 => n5221, C2 => 
                           MEM_IN(9), A => n5264_port, ZN => n5263_port);
   U5704 : OAI22_X1 port map( A1 => n11748, A2 => n231, B1 => n4961, B2 => 
                           n5224, ZN => n5264_port);
   U5705 : AOI22_X1 port map( A1 => n5225, A2 => n4962, B1 => n5226, B2 => 
                           n4963, ZN => n5262_port);
   U5706 : AOI22_X1 port map( A1 => n5227, A2 => n4964, B1 => n5228, B2 => 
                           n4965, ZN => n5261_port);
   U5707 : NAND3_X1 port map( A1 => n5265_port, A2 => n5266_port, A3 => 
                           n5267_port, ZN => n13110);
   U5708 : AOI221_X1 port map( B1 => n5220, B2 => n4969, C1 => n5221, C2 => 
                           MEM_IN(10), A => n5268_port, ZN => n5267_port);
   U5709 : OAI22_X1 port map( A1 => n11747, A2 => n231, B1 => n4971, B2 => 
                           n5224, ZN => n5268_port);
   U5710 : AOI22_X1 port map( A1 => n5225, A2 => n4972, B1 => n5226, B2 => 
                           n4973, ZN => n5266_port);
   U5711 : AOI22_X1 port map( A1 => n5227, A2 => n4974, B1 => n5228, B2 => 
                           n4975, ZN => n5265_port);
   U5712 : NAND3_X1 port map( A1 => n5269_port, A2 => n5270_port, A3 => 
                           n5271_port, ZN => n13109);
   U5713 : AOI221_X1 port map( B1 => n5220, B2 => n4979, C1 => n5221, C2 => 
                           MEM_IN(11), A => n5272_port, ZN => n5271_port);
   U5714 : OAI22_X1 port map( A1 => n11746, A2 => n231, B1 => n4981, B2 => 
                           n5224, ZN => n5272_port);
   U5715 : AOI22_X1 port map( A1 => n5225, A2 => n4982, B1 => n5226, B2 => 
                           n4983, ZN => n5270_port);
   U5716 : AOI22_X1 port map( A1 => n5227, A2 => n4984, B1 => n5228, B2 => 
                           n4985, ZN => n5269_port);
   U5717 : NAND3_X1 port map( A1 => n5273_port, A2 => n5274_port, A3 => 
                           n5275_port, ZN => n13108);
   U5718 : AOI221_X1 port map( B1 => n5220, B2 => n4989, C1 => n5221, C2 => 
                           MEM_IN(12), A => n5276_port, ZN => n5275_port);
   U5719 : OAI22_X1 port map( A1 => n11745, A2 => n231, B1 => n4991, B2 => 
                           n5224, ZN => n5276_port);
   U5720 : AOI22_X1 port map( A1 => n5225, A2 => n4992, B1 => n5226, B2 => 
                           n4993, ZN => n5274_port);
   U5721 : AOI22_X1 port map( A1 => n5227, A2 => n4994, B1 => n5228, B2 => 
                           n4995, ZN => n5273_port);
   U5722 : NAND3_X1 port map( A1 => n5277_port, A2 => n5278_port, A3 => 
                           n5279_port, ZN => n13107);
   U5723 : AOI221_X1 port map( B1 => n5220, B2 => n4999, C1 => n5221, C2 => 
                           MEM_IN(13), A => n5280_port, ZN => n5279_port);
   U5724 : OAI22_X1 port map( A1 => n11744, A2 => n231, B1 => n5001, B2 => 
                           n5224, ZN => n5280_port);
   U5725 : AOI22_X1 port map( A1 => n5225, A2 => n5002, B1 => n5226, B2 => 
                           n5003, ZN => n5278_port);
   U5726 : AOI22_X1 port map( A1 => n5227, A2 => n5004, B1 => n5228, B2 => 
                           n5005, ZN => n5277_port);
   U5727 : NAND3_X1 port map( A1 => n5281_port, A2 => n5282, A3 => n5283, ZN =>
                           n13106);
   U5728 : AOI221_X1 port map( B1 => n5220, B2 => n5009, C1 => n5221, C2 => 
                           MEM_IN(14), A => n5284, ZN => n5283);
   U5729 : OAI22_X1 port map( A1 => n11743, A2 => n231, B1 => n5011, B2 => 
                           n5224, ZN => n5284);
   U5730 : AOI22_X1 port map( A1 => n5225, A2 => n5012, B1 => n5226, B2 => 
                           n5013, ZN => n5282);
   U5731 : AOI22_X1 port map( A1 => n5227, A2 => n5014, B1 => n5228, B2 => 
                           n5015, ZN => n5281_port);
   U5732 : NAND3_X1 port map( A1 => n5285, A2 => n5286, A3 => n5287, ZN => 
                           n13105);
   U5733 : AOI221_X1 port map( B1 => n5220, B2 => n5019, C1 => n5221, C2 => 
                           MEM_IN(15), A => n5288, ZN => n5287);
   U5734 : OAI22_X1 port map( A1 => n11742, A2 => n231, B1 => n5021, B2 => 
                           n5224, ZN => n5288);
   U5735 : AOI22_X1 port map( A1 => n5225, A2 => n5022, B1 => n5226, B2 => 
                           n5023, ZN => n5286);
   U5736 : AOI22_X1 port map( A1 => n5227, A2 => n5024, B1 => n5228, B2 => 
                           n5025, ZN => n5285);
   U5737 : NAND3_X1 port map( A1 => n5289, A2 => n5290, A3 => n5291, ZN => 
                           n13104);
   U5738 : AOI221_X1 port map( B1 => n5220, B2 => n5029, C1 => n5221, C2 => 
                           MEM_IN(16), A => n5292, ZN => n5291);
   U5739 : OAI22_X1 port map( A1 => n11741, A2 => n231, B1 => n5031, B2 => 
                           n5224, ZN => n5292);
   U5740 : AOI22_X1 port map( A1 => n5225, A2 => n5032, B1 => n5226, B2 => 
                           n5033, ZN => n5290);
   U5741 : AOI22_X1 port map( A1 => n5227, A2 => n5034, B1 => n5228, B2 => 
                           n5035, ZN => n5289);
   U5742 : NAND3_X1 port map( A1 => n5293, A2 => n5294, A3 => n5295, ZN => 
                           n13103);
   U5743 : AOI221_X1 port map( B1 => n5220, B2 => n5039, C1 => n5221, C2 => 
                           MEM_IN(17), A => n5296, ZN => n5295);
   U5744 : OAI22_X1 port map( A1 => n11740, A2 => n231, B1 => n5041, B2 => 
                           n5224, ZN => n5296);
   U5745 : AOI22_X1 port map( A1 => n5225, A2 => n5042, B1 => n5226, B2 => 
                           n5043, ZN => n5294);
   U5746 : AOI22_X1 port map( A1 => n5227, A2 => n5044, B1 => n5228, B2 => 
                           n5045, ZN => n5293);
   U5747 : NAND3_X1 port map( A1 => n5297, A2 => n5298, A3 => n5299, ZN => 
                           n13102);
   U5748 : AOI221_X1 port map( B1 => n5220, B2 => n5049, C1 => n5221, C2 => 
                           MEM_IN(18), A => n5300, ZN => n5299);
   U5749 : OAI22_X1 port map( A1 => n11739, A2 => n231, B1 => n5051, B2 => 
                           n5224, ZN => n5300);
   U5750 : AOI22_X1 port map( A1 => n5225, A2 => n5052, B1 => n5226, B2 => 
                           n5053, ZN => n5298);
   U5751 : AOI22_X1 port map( A1 => n5227, A2 => n5054, B1 => n5228, B2 => 
                           n5055, ZN => n5297);
   U5752 : NAND3_X1 port map( A1 => n5301, A2 => n5302, A3 => n5303, ZN => 
                           n13101);
   U5753 : AOI221_X1 port map( B1 => n5220, B2 => n5059, C1 => n5221, C2 => 
                           MEM_IN(19), A => n5304, ZN => n5303);
   U5754 : OAI22_X1 port map( A1 => n11738, A2 => n231, B1 => n5061, B2 => 
                           n5224, ZN => n5304);
   U5755 : AOI22_X1 port map( A1 => n5225, A2 => n5062, B1 => n5226, B2 => 
                           n5063, ZN => n5302);
   U5756 : AOI22_X1 port map( A1 => n5227, A2 => n5064, B1 => n5228, B2 => 
                           n5065, ZN => n5301);
   U5757 : NAND3_X1 port map( A1 => n5305, A2 => n5306, A3 => n5307, ZN => 
                           n13100);
   U5758 : AOI221_X1 port map( B1 => n5220, B2 => n5069, C1 => n5221, C2 => 
                           MEM_IN(20), A => n5308, ZN => n5307);
   U5759 : OAI22_X1 port map( A1 => n11737, A2 => n231, B1 => n5071, B2 => 
                           n5224, ZN => n5308);
   U5760 : AOI22_X1 port map( A1 => n5225, A2 => n5072, B1 => n5226, B2 => 
                           n5073, ZN => n5306);
   U5761 : AOI22_X1 port map( A1 => n5227, A2 => n5074, B1 => n5228, B2 => 
                           n5075, ZN => n5305);
   U5762 : NAND3_X1 port map( A1 => n5309, A2 => n5310, A3 => n5311, ZN => 
                           n13099);
   U5763 : AOI221_X1 port map( B1 => n5220, B2 => n5079, C1 => n5221, C2 => 
                           MEM_IN(21), A => n5312, ZN => n5311);
   U5764 : OAI22_X1 port map( A1 => n11736, A2 => n231, B1 => n5081, B2 => 
                           n5224, ZN => n5312);
   U5765 : AOI22_X1 port map( A1 => n5225, A2 => n5082, B1 => n5226, B2 => 
                           n5083, ZN => n5310);
   U5766 : AOI22_X1 port map( A1 => n5227, A2 => n5084, B1 => n5228, B2 => 
                           n5085, ZN => n5309);
   U5767 : NAND3_X1 port map( A1 => n5313, A2 => n5314, A3 => n5315, ZN => 
                           n13098);
   U5768 : AOI221_X1 port map( B1 => n5220, B2 => n5089, C1 => n5221, C2 => 
                           MEM_IN(22), A => n5316, ZN => n5315);
   U5769 : OAI22_X1 port map( A1 => n11735, A2 => n231, B1 => n5091, B2 => 
                           n5224, ZN => n5316);
   U5770 : AOI22_X1 port map( A1 => n5225, A2 => n5092, B1 => n5226, B2 => 
                           n5093, ZN => n5314);
   U5771 : AOI22_X1 port map( A1 => n5227, A2 => n5094, B1 => n5228, B2 => 
                           n5095, ZN => n5313);
   U5772 : NAND3_X1 port map( A1 => n5317, A2 => n5318, A3 => n5319, ZN => 
                           n13097);
   U5773 : AOI221_X1 port map( B1 => n5220, B2 => n5099, C1 => n5221, C2 => 
                           MEM_IN(23), A => n5320, ZN => n5319);
   U5774 : OAI22_X1 port map( A1 => n11734, A2 => n231, B1 => n5101, B2 => 
                           n5224, ZN => n5320);
   U5775 : AOI22_X1 port map( A1 => n5225, A2 => n5102, B1 => n5226, B2 => 
                           n5103, ZN => n5318);
   U5776 : AOI22_X1 port map( A1 => n5227, A2 => n5104, B1 => n5228, B2 => 
                           n5105, ZN => n5317);
   U5777 : NAND3_X1 port map( A1 => n5321, A2 => n5322, A3 => n5323, ZN => 
                           n13096);
   U5778 : AOI221_X1 port map( B1 => n5220, B2 => n5109, C1 => n5221, C2 => 
                           MEM_IN(24), A => n5324, ZN => n5323);
   U5779 : OAI22_X1 port map( A1 => n11733, A2 => n231, B1 => n5111, B2 => 
                           n5224, ZN => n5324);
   U5780 : AOI22_X1 port map( A1 => n5225, A2 => n5112, B1 => n5226, B2 => 
                           n5113, ZN => n5322);
   U5781 : AOI22_X1 port map( A1 => n5227, A2 => n5114, B1 => n5228, B2 => 
                           n5115, ZN => n5321);
   U5782 : NAND3_X1 port map( A1 => n5325, A2 => n5326, A3 => n5327, ZN => 
                           n13095);
   U5783 : AOI221_X1 port map( B1 => n5220, B2 => n5119, C1 => n5221, C2 => 
                           MEM_IN(25), A => n5328, ZN => n5327);
   U5784 : OAI22_X1 port map( A1 => n11732, A2 => n231, B1 => n5121, B2 => 
                           n5224, ZN => n5328);
   U5785 : AOI22_X1 port map( A1 => n5225, A2 => n5122, B1 => n5226, B2 => 
                           n5123, ZN => n5326);
   U5786 : AOI22_X1 port map( A1 => n5227, A2 => n5124, B1 => n5228, B2 => 
                           n5125, ZN => n5325);
   U5787 : NAND3_X1 port map( A1 => n5329, A2 => n5330, A3 => n5331, ZN => 
                           n13094);
   U5788 : AOI221_X1 port map( B1 => n5220, B2 => n5129, C1 => n5221, C2 => 
                           MEM_IN(26), A => n5332, ZN => n5331);
   U5789 : OAI22_X1 port map( A1 => n11731, A2 => n231, B1 => n5131, B2 => 
                           n5224, ZN => n5332);
   U5790 : AOI22_X1 port map( A1 => n5225, A2 => n5132, B1 => n5226, B2 => 
                           n5133, ZN => n5330);
   U5791 : AOI22_X1 port map( A1 => n5227, A2 => n5134, B1 => n5228, B2 => 
                           n5135, ZN => n5329);
   U5792 : NAND3_X1 port map( A1 => n5333, A2 => n5334, A3 => n5335, ZN => 
                           n13093);
   U5793 : AOI221_X1 port map( B1 => n5220, B2 => n5139, C1 => n5221, C2 => 
                           MEM_IN(27), A => n5336, ZN => n5335);
   U5794 : OAI22_X1 port map( A1 => n11730, A2 => n231, B1 => n5141, B2 => 
                           n5224, ZN => n5336);
   U5795 : AOI22_X1 port map( A1 => n5225, A2 => n5142, B1 => n5226, B2 => 
                           n5143, ZN => n5334);
   U5796 : AOI22_X1 port map( A1 => n5227, A2 => n5144, B1 => n5228, B2 => 
                           n5145, ZN => n5333);
   U5797 : NAND3_X1 port map( A1 => n5337, A2 => n5338, A3 => n5339, ZN => 
                           n13092);
   U5798 : AOI221_X1 port map( B1 => n5220, B2 => n5149, C1 => n5221, C2 => 
                           MEM_IN(28), A => n5340, ZN => n5339);
   U5799 : OAI22_X1 port map( A1 => n11729, A2 => n231, B1 => n5151, B2 => 
                           n5224, ZN => n5340);
   U5800 : AOI22_X1 port map( A1 => n5225, A2 => n5152, B1 => n5226, B2 => 
                           n5153, ZN => n5338);
   U5801 : AOI22_X1 port map( A1 => n5227, A2 => n5154, B1 => n5228, B2 => 
                           n5155, ZN => n5337);
   U5802 : NAND3_X1 port map( A1 => n5341, A2 => n5342, A3 => n5343, ZN => 
                           n13091);
   U5803 : AOI221_X1 port map( B1 => n5220, B2 => n5159, C1 => n5221, C2 => 
                           MEM_IN(29), A => n5344, ZN => n5343);
   U5804 : OAI22_X1 port map( A1 => n11728, A2 => n231, B1 => n5161, B2 => 
                           n5224, ZN => n5344);
   U5805 : AOI22_X1 port map( A1 => n5225, A2 => n5162, B1 => n5226, B2 => 
                           n5163, ZN => n5342);
   U5806 : AOI22_X1 port map( A1 => n5227, A2 => n5164, B1 => n5228, B2 => 
                           n5165, ZN => n5341);
   U5807 : NAND3_X1 port map( A1 => n5345, A2 => n5346, A3 => n5347, ZN => 
                           n13090);
   U5808 : AOI221_X1 port map( B1 => n5220, B2 => n5169, C1 => n5221, C2 => 
                           MEM_IN(30), A => n5348, ZN => n5347);
   U5809 : OAI22_X1 port map( A1 => n11727, A2 => n231, B1 => n5171, B2 => 
                           n5224, ZN => n5348);
   U5810 : AOI22_X1 port map( A1 => n5225, A2 => n5172, B1 => n5226, B2 => 
                           n5173, ZN => n5346);
   U5811 : AOI22_X1 port map( A1 => n5227, A2 => n5174, B1 => n5228, B2 => 
                           n5175, ZN => n5345);
   U5812 : NAND3_X1 port map( A1 => n5349, A2 => n5350, A3 => n5351, ZN => 
                           n13089);
   U5813 : AOI221_X1 port map( B1 => n5220, B2 => n5179, C1 => n5221, C2 => 
                           MEM_IN(31), A => n5352, ZN => n5351);
   U5814 : OAI22_X1 port map( A1 => n11726, A2 => n231, B1 => n5181, B2 => 
                           n5224, ZN => n5352);
   U5815 : OAI21_X1 port map( B1 => n5357, B2 => n4787, A => n5358, ZN => n5356
                           );
   U5816 : NOR3_X1 port map( A1 => n5188, A2 => n5359, A3 => n5190, ZN => n5357
                           );
   U5817 : AOI22_X1 port map( A1 => n5225, A2 => n5191, B1 => n5226, B2 => 
                           n5192, ZN => n5350);
   U5818 : AOI22_X1 port map( A1 => n5227, A2 => n5195, B1 => n5228, B2 => 
                           n5196, ZN => n5349);
   U5819 : OAI22_X1 port map( A1 => n5355, A2 => n5361, B1 => n208, B2 => n230,
                           ZN => n5358);
   U5820 : INV_X1 port map( A => n5354, ZN => n5361);
   U5821 : NOR3_X1 port map( A1 => n4841, A2 => n230, A3 => n5353, ZN => n5354)
                           ;
   U5822 : OAI22_X1 port map( A1 => n4786, A2 => n5362, B1 => n5363, B2 => 
                           n5204, ZN => n5223);
   U5823 : NOR2_X1 port map( A1 => n5353, A2 => n5355, ZN => n5363);
   U5824 : NAND2_X1 port map( A1 => n5364, A2 => n5212, ZN => n5353);
   U5825 : AOI211_X1 port map( C1 => n5208, C2 => n5365, A => n5209, B => n5360
                           , ZN => n5362);
   U5826 : OAI211_X1 port map( C1 => n5366, C2 => n4787, A => n5367, B => n5368
                           , ZN => n5209);
   U5827 : INV_X1 port map( A => n5188, ZN => n5366);
   U5828 : NAND2_X1 port map( A1 => n5369, A2 => n5212, ZN => n5188);
   U5829 : OR2_X1 port map( A1 => n5370, A2 => n5371, ZN => n5355);
   U5830 : NOR2_X1 port map( A1 => n5212, A2 => n5190, ZN => n5197);
   U5831 : NAND2_X1 port map( A1 => n5372, A2 => n5216, ZN => n5212);
   U5832 : NAND3_X1 port map( A1 => n5373, A2 => n5374, A3 => n5375, ZN => 
                           n13088);
   U5833 : AOI221_X1 port map( B1 => n5376, B2 => n4863, C1 => n5377, C2 => 
                           MEM_IN(0), A => n5378, ZN => n5375);
   U5834 : OAI22_X1 port map( A1 => n11725, A2 => n233, B1 => n4867, B2 => 
                           n5380, ZN => n5378);
   U5835 : AOI22_X1 port map( A1 => n5381, A2 => n4869, B1 => n5382, B2 => 
                           n4871, ZN => n5374);
   U5836 : AOI22_X1 port map( A1 => n5383, A2 => n4873, B1 => n5384, B2 => 
                           n4875, ZN => n5373);
   U5837 : NAND3_X1 port map( A1 => n5385, A2 => n5386, A3 => n5387, ZN => 
                           n13087);
   U5838 : AOI221_X1 port map( B1 => n5376, B2 => n4879, C1 => n5377, C2 => 
                           MEM_IN(1), A => n5388, ZN => n5387);
   U5839 : OAI22_X1 port map( A1 => n11724, A2 => n233, B1 => n4881, B2 => 
                           n5380, ZN => n5388);
   U5840 : AOI22_X1 port map( A1 => n5381, A2 => n4882, B1 => n5382, B2 => 
                           n4883, ZN => n5386);
   U5841 : AOI22_X1 port map( A1 => n5383, A2 => n4884, B1 => n5384, B2 => 
                           n4885, ZN => n5385);
   U5842 : NAND3_X1 port map( A1 => n5389, A2 => n5390, A3 => n5391, ZN => 
                           n13086);
   U5843 : AOI221_X1 port map( B1 => n5376, B2 => n4889, C1 => n5377, C2 => 
                           MEM_IN(2), A => n5392, ZN => n5391);
   U5844 : OAI22_X1 port map( A1 => n11723, A2 => n233, B1 => n4891, B2 => 
                           n5380, ZN => n5392);
   U5845 : AOI22_X1 port map( A1 => n5381, A2 => n4892, B1 => n5382, B2 => 
                           n4893, ZN => n5390);
   U5846 : AOI22_X1 port map( A1 => n5383, A2 => n4894, B1 => n5384, B2 => 
                           n4895, ZN => n5389);
   U5847 : NAND3_X1 port map( A1 => n5393, A2 => n5394, A3 => n5395, ZN => 
                           n13085);
   U5848 : AOI221_X1 port map( B1 => n5376, B2 => n4899, C1 => n5377, C2 => 
                           MEM_IN(3), A => n5396, ZN => n5395);
   U5849 : OAI22_X1 port map( A1 => n11722, A2 => n233, B1 => n4901, B2 => 
                           n5380, ZN => n5396);
   U5850 : AOI22_X1 port map( A1 => n5381, A2 => n4902, B1 => n5382, B2 => 
                           n4903, ZN => n5394);
   U5851 : AOI22_X1 port map( A1 => n5383, A2 => n4904, B1 => n5384, B2 => 
                           n4905, ZN => n5393);
   U5852 : NAND3_X1 port map( A1 => n5397, A2 => n5398, A3 => n5399, ZN => 
                           n13084);
   U5853 : AOI221_X1 port map( B1 => n5376, B2 => n4909, C1 => n5377, C2 => 
                           MEM_IN(4), A => n5400, ZN => n5399);
   U5854 : OAI22_X1 port map( A1 => n11721, A2 => n233, B1 => n4911, B2 => 
                           n5380, ZN => n5400);
   U5855 : AOI22_X1 port map( A1 => n5381, A2 => n4912, B1 => n5382, B2 => 
                           n4913, ZN => n5398);
   U5856 : AOI22_X1 port map( A1 => n5383, A2 => n4914, B1 => n5384, B2 => 
                           n4915, ZN => n5397);
   U5857 : NAND3_X1 port map( A1 => n5401, A2 => n5402, A3 => n5403, ZN => 
                           n13083);
   U5858 : AOI221_X1 port map( B1 => n5376, B2 => n4919, C1 => n5377, C2 => 
                           MEM_IN(5), A => n5404, ZN => n5403);
   U5859 : OAI22_X1 port map( A1 => n11720, A2 => n233, B1 => n4921, B2 => 
                           n5380, ZN => n5404);
   U5860 : AOI22_X1 port map( A1 => n5381, A2 => n4922, B1 => n5382, B2 => 
                           n4923, ZN => n5402);
   U5861 : AOI22_X1 port map( A1 => n5383, A2 => n4924, B1 => n5384, B2 => 
                           n4925, ZN => n5401);
   U5862 : NAND3_X1 port map( A1 => n5405, A2 => n5406, A3 => n5407, ZN => 
                           n13082);
   U5863 : AOI221_X1 port map( B1 => n5376, B2 => n4929, C1 => n5377, C2 => 
                           MEM_IN(6), A => n5408, ZN => n5407);
   U5864 : OAI22_X1 port map( A1 => n11719, A2 => n233, B1 => n4931, B2 => 
                           n5380, ZN => n5408);
   U5865 : AOI22_X1 port map( A1 => n5381, A2 => n4932, B1 => n5382, B2 => 
                           n4933, ZN => n5406);
   U5866 : AOI22_X1 port map( A1 => n5383, A2 => n4934, B1 => n5384, B2 => 
                           n4935, ZN => n5405);
   U5867 : NAND3_X1 port map( A1 => n5409, A2 => n5410, A3 => n5411, ZN => 
                           n13081);
   U5868 : AOI221_X1 port map( B1 => n5376, B2 => n4939, C1 => n5377, C2 => 
                           MEM_IN(7), A => n5412, ZN => n5411);
   U5869 : OAI22_X1 port map( A1 => n11718, A2 => n233, B1 => n4941, B2 => 
                           n5380, ZN => n5412);
   U5870 : AOI22_X1 port map( A1 => n5381, A2 => n4942, B1 => n5382, B2 => 
                           n4943, ZN => n5410);
   U5871 : AOI22_X1 port map( A1 => n5383, A2 => n4944, B1 => n5384, B2 => 
                           n4945, ZN => n5409);
   U5872 : NAND3_X1 port map( A1 => n5413, A2 => n5414, A3 => n5415, ZN => 
                           n13080);
   U5873 : AOI221_X1 port map( B1 => n5376, B2 => n4949, C1 => n5377, C2 => 
                           MEM_IN(8), A => n5416, ZN => n5415);
   U5874 : OAI22_X1 port map( A1 => n11717, A2 => n233, B1 => n4951, B2 => 
                           n5380, ZN => n5416);
   U5875 : AOI22_X1 port map( A1 => n5381, A2 => n4952, B1 => n5382, B2 => 
                           n4953, ZN => n5414);
   U5876 : AOI22_X1 port map( A1 => n5383, A2 => n4954, B1 => n5384, B2 => 
                           n4955, ZN => n5413);
   U5877 : NAND3_X1 port map( A1 => n5417, A2 => n5418, A3 => n5419, ZN => 
                           n13079);
   U5878 : AOI221_X1 port map( B1 => n5376, B2 => n4959, C1 => n5377, C2 => 
                           MEM_IN(9), A => n5420, ZN => n5419);
   U5879 : OAI22_X1 port map( A1 => n11716, A2 => n233, B1 => n4961, B2 => 
                           n5380, ZN => n5420);
   U5880 : AOI22_X1 port map( A1 => n5381, A2 => n4962, B1 => n5382, B2 => 
                           n4963, ZN => n5418);
   U5881 : AOI22_X1 port map( A1 => n5383, A2 => n4964, B1 => n5384, B2 => 
                           n4965, ZN => n5417);
   U5882 : NAND3_X1 port map( A1 => n5421, A2 => n5422, A3 => n5423, ZN => 
                           n13078);
   U5883 : AOI221_X1 port map( B1 => n5376, B2 => n4969, C1 => n5377, C2 => 
                           MEM_IN(10), A => n5424, ZN => n5423);
   U5884 : OAI22_X1 port map( A1 => n11715, A2 => n233, B1 => n4971, B2 => 
                           n5380, ZN => n5424);
   U5885 : AOI22_X1 port map( A1 => n5381, A2 => n4972, B1 => n5382, B2 => 
                           n4973, ZN => n5422);
   U5886 : AOI22_X1 port map( A1 => n5383, A2 => n4974, B1 => n5384, B2 => 
                           n4975, ZN => n5421);
   U5887 : NAND3_X1 port map( A1 => n5425, A2 => n5426, A3 => n5427, ZN => 
                           n13077);
   U5888 : AOI221_X1 port map( B1 => n5376, B2 => n4979, C1 => n5377, C2 => 
                           MEM_IN(11), A => n5428, ZN => n5427);
   U5889 : OAI22_X1 port map( A1 => n11714, A2 => n233, B1 => n4981, B2 => 
                           n5380, ZN => n5428);
   U5890 : AOI22_X1 port map( A1 => n5381, A2 => n4982, B1 => n5382, B2 => 
                           n4983, ZN => n5426);
   U5891 : AOI22_X1 port map( A1 => n5383, A2 => n4984, B1 => n5384, B2 => 
                           n4985, ZN => n5425);
   U5892 : NAND3_X1 port map( A1 => n5429, A2 => n5430, A3 => n5431, ZN => 
                           n13076);
   U5893 : AOI221_X1 port map( B1 => n5376, B2 => n4989, C1 => n5377, C2 => 
                           MEM_IN(12), A => n5432, ZN => n5431);
   U5894 : OAI22_X1 port map( A1 => n11713, A2 => n233, B1 => n4991, B2 => 
                           n5380, ZN => n5432);
   U5895 : AOI22_X1 port map( A1 => n5381, A2 => n4992, B1 => n5382, B2 => 
                           n4993, ZN => n5430);
   U5896 : AOI22_X1 port map( A1 => n5383, A2 => n4994, B1 => n5384, B2 => 
                           n4995, ZN => n5429);
   U5897 : NAND3_X1 port map( A1 => n5433, A2 => n5434, A3 => n5435, ZN => 
                           n13075);
   U5898 : AOI221_X1 port map( B1 => n5376, B2 => n4999, C1 => n5377, C2 => 
                           MEM_IN(13), A => n5436, ZN => n5435);
   U5899 : OAI22_X1 port map( A1 => n11712, A2 => n233, B1 => n5001, B2 => 
                           n5380, ZN => n5436);
   U5900 : AOI22_X1 port map( A1 => n5381, A2 => n5002, B1 => n5382, B2 => 
                           n5003, ZN => n5434);
   U5901 : AOI22_X1 port map( A1 => n5383, A2 => n5004, B1 => n5384, B2 => 
                           n5005, ZN => n5433);
   U5902 : NAND3_X1 port map( A1 => n5437, A2 => n5438, A3 => n5439, ZN => 
                           n13074);
   U5903 : AOI221_X1 port map( B1 => n5376, B2 => n5009, C1 => n5377, C2 => 
                           MEM_IN(14), A => n5440, ZN => n5439);
   U5904 : OAI22_X1 port map( A1 => n11711, A2 => n233, B1 => n5011, B2 => 
                           n5380, ZN => n5440);
   U5905 : AOI22_X1 port map( A1 => n5381, A2 => n5012, B1 => n5382, B2 => 
                           n5013, ZN => n5438);
   U5906 : AOI22_X1 port map( A1 => n5383, A2 => n5014, B1 => n5384, B2 => 
                           n5015, ZN => n5437);
   U5907 : NAND3_X1 port map( A1 => n5441, A2 => n5442, A3 => n5443, ZN => 
                           n13073);
   U5908 : AOI221_X1 port map( B1 => n5376, B2 => n5019, C1 => n5377, C2 => 
                           MEM_IN(15), A => n5444, ZN => n5443);
   U5909 : OAI22_X1 port map( A1 => n11710, A2 => n233, B1 => n5021, B2 => 
                           n5380, ZN => n5444);
   U5910 : AOI22_X1 port map( A1 => n5381, A2 => n5022, B1 => n5382, B2 => 
                           n5023, ZN => n5442);
   U5911 : AOI22_X1 port map( A1 => n5383, A2 => n5024, B1 => n5384, B2 => 
                           n5025, ZN => n5441);
   U5912 : NAND3_X1 port map( A1 => n5445, A2 => n5446, A3 => n5447, ZN => 
                           n13072);
   U5913 : AOI221_X1 port map( B1 => n5376, B2 => n5029, C1 => n5377, C2 => 
                           MEM_IN(16), A => n5448, ZN => n5447);
   U5914 : OAI22_X1 port map( A1 => n11709, A2 => n233, B1 => n5031, B2 => 
                           n5380, ZN => n5448);
   U5915 : AOI22_X1 port map( A1 => n5381, A2 => n5032, B1 => n5382, B2 => 
                           n5033, ZN => n5446);
   U5916 : AOI22_X1 port map( A1 => n5383, A2 => n5034, B1 => n5384, B2 => 
                           n5035, ZN => n5445);
   U5917 : NAND3_X1 port map( A1 => n5449, A2 => n5450, A3 => n5451, ZN => 
                           n13071);
   U5918 : AOI221_X1 port map( B1 => n5376, B2 => n5039, C1 => n5377, C2 => 
                           MEM_IN(17), A => n5452, ZN => n5451);
   U5919 : OAI22_X1 port map( A1 => n11708, A2 => n233, B1 => n5041, B2 => 
                           n5380, ZN => n5452);
   U5920 : AOI22_X1 port map( A1 => n5381, A2 => n5042, B1 => n5382, B2 => 
                           n5043, ZN => n5450);
   U5921 : AOI22_X1 port map( A1 => n5383, A2 => n5044, B1 => n5384, B2 => 
                           n5045, ZN => n5449);
   U5922 : NAND3_X1 port map( A1 => n5453, A2 => n5454, A3 => n5455, ZN => 
                           n13070);
   U5923 : AOI221_X1 port map( B1 => n5376, B2 => n5049, C1 => n5377, C2 => 
                           MEM_IN(18), A => n5456, ZN => n5455);
   U5924 : OAI22_X1 port map( A1 => n11707, A2 => n233, B1 => n5051, B2 => 
                           n5380, ZN => n5456);
   U5925 : AOI22_X1 port map( A1 => n5381, A2 => n5052, B1 => n5382, B2 => 
                           n5053, ZN => n5454);
   U5926 : AOI22_X1 port map( A1 => n5383, A2 => n5054, B1 => n5384, B2 => 
                           n5055, ZN => n5453);
   U5927 : NAND3_X1 port map( A1 => n5457, A2 => n5458, A3 => n5459, ZN => 
                           n13069);
   U5928 : AOI221_X1 port map( B1 => n5376, B2 => n5059, C1 => n5377, C2 => 
                           MEM_IN(19), A => n5460, ZN => n5459);
   U5929 : OAI22_X1 port map( A1 => n11706, A2 => n233, B1 => n5061, B2 => 
                           n5380, ZN => n5460);
   U5930 : AOI22_X1 port map( A1 => n5381, A2 => n5062, B1 => n5382, B2 => 
                           n5063, ZN => n5458);
   U5931 : AOI22_X1 port map( A1 => n5383, A2 => n5064, B1 => n5384, B2 => 
                           n5065, ZN => n5457);
   U5932 : NAND3_X1 port map( A1 => n5461, A2 => n5462, A3 => n5463, ZN => 
                           n13068);
   U5933 : AOI221_X1 port map( B1 => n5376, B2 => n5069, C1 => n5377, C2 => 
                           MEM_IN(20), A => n5464, ZN => n5463);
   U5934 : OAI22_X1 port map( A1 => n11705, A2 => n233, B1 => n5071, B2 => 
                           n5380, ZN => n5464);
   U5935 : AOI22_X1 port map( A1 => n5381, A2 => n5072, B1 => n5382, B2 => 
                           n5073, ZN => n5462);
   U5936 : AOI22_X1 port map( A1 => n5383, A2 => n5074, B1 => n5384, B2 => 
                           n5075, ZN => n5461);
   U5937 : NAND3_X1 port map( A1 => n5465, A2 => n5466, A3 => n5467, ZN => 
                           n13067);
   U5938 : AOI221_X1 port map( B1 => n5376, B2 => n5079, C1 => n5377, C2 => 
                           MEM_IN(21), A => n5468, ZN => n5467);
   U5939 : OAI22_X1 port map( A1 => n11704, A2 => n233, B1 => n5081, B2 => 
                           n5380, ZN => n5468);
   U5940 : AOI22_X1 port map( A1 => n5381, A2 => n5082, B1 => n5382, B2 => 
                           n5083, ZN => n5466);
   U5941 : AOI22_X1 port map( A1 => n5383, A2 => n5084, B1 => n5384, B2 => 
                           n5085, ZN => n5465);
   U5942 : NAND3_X1 port map( A1 => n5469, A2 => n5470, A3 => n5471, ZN => 
                           n13066);
   U5943 : AOI221_X1 port map( B1 => n5376, B2 => n5089, C1 => n5377, C2 => 
                           MEM_IN(22), A => n5472, ZN => n5471);
   U5944 : OAI22_X1 port map( A1 => n11703, A2 => n233, B1 => n5091, B2 => 
                           n5380, ZN => n5472);
   U5945 : AOI22_X1 port map( A1 => n5381, A2 => n5092, B1 => n5382, B2 => 
                           n5093, ZN => n5470);
   U5946 : AOI22_X1 port map( A1 => n5383, A2 => n5094, B1 => n5384, B2 => 
                           n5095, ZN => n5469);
   U5947 : NAND3_X1 port map( A1 => n5473, A2 => n5474, A3 => n5475, ZN => 
                           n13065);
   U5948 : AOI221_X1 port map( B1 => n5376, B2 => n5099, C1 => n5377, C2 => 
                           MEM_IN(23), A => n5476, ZN => n5475);
   U5949 : OAI22_X1 port map( A1 => n11702, A2 => n233, B1 => n5101, B2 => 
                           n5380, ZN => n5476);
   U5950 : AOI22_X1 port map( A1 => n5381, A2 => n5102, B1 => n5382, B2 => 
                           n5103, ZN => n5474);
   U5951 : AOI22_X1 port map( A1 => n5383, A2 => n5104, B1 => n5384, B2 => 
                           n5105, ZN => n5473);
   U5952 : NAND3_X1 port map( A1 => n5477, A2 => n5478, A3 => n5479, ZN => 
                           n13064);
   U5953 : AOI221_X1 port map( B1 => n5376, B2 => n5109, C1 => n5377, C2 => 
                           MEM_IN(24), A => n5480, ZN => n5479);
   U5954 : OAI22_X1 port map( A1 => n11701, A2 => n233, B1 => n5111, B2 => 
                           n5380, ZN => n5480);
   U5955 : AOI22_X1 port map( A1 => n5381, A2 => n5112, B1 => n5382, B2 => 
                           n5113, ZN => n5478);
   U5956 : AOI22_X1 port map( A1 => n5383, A2 => n5114, B1 => n5384, B2 => 
                           n5115, ZN => n5477);
   U5957 : NAND3_X1 port map( A1 => n5481, A2 => n5482, A3 => n5483, ZN => 
                           n13063);
   U5958 : AOI221_X1 port map( B1 => n5376, B2 => n5119, C1 => n5377, C2 => 
                           MEM_IN(25), A => n5484, ZN => n5483);
   U5959 : OAI22_X1 port map( A1 => n11700, A2 => n233, B1 => n5121, B2 => 
                           n5380, ZN => n5484);
   U5960 : AOI22_X1 port map( A1 => n5381, A2 => n5122, B1 => n5382, B2 => 
                           n5123, ZN => n5482);
   U5961 : AOI22_X1 port map( A1 => n5383, A2 => n5124, B1 => n5384, B2 => 
                           n5125, ZN => n5481);
   U5962 : NAND3_X1 port map( A1 => n5485, A2 => n5486, A3 => n5487, ZN => 
                           n13062);
   U5963 : AOI221_X1 port map( B1 => n5376, B2 => n5129, C1 => n5377, C2 => 
                           MEM_IN(26), A => n5488, ZN => n5487);
   U5964 : OAI22_X1 port map( A1 => n11699, A2 => n233, B1 => n5131, B2 => 
                           n5380, ZN => n5488);
   U5965 : AOI22_X1 port map( A1 => n5381, A2 => n5132, B1 => n5382, B2 => 
                           n5133, ZN => n5486);
   U5966 : AOI22_X1 port map( A1 => n5383, A2 => n5134, B1 => n5384, B2 => 
                           n5135, ZN => n5485);
   U5967 : NAND3_X1 port map( A1 => n5489, A2 => n5490, A3 => n5491, ZN => 
                           n13061);
   U5968 : AOI221_X1 port map( B1 => n5376, B2 => n5139, C1 => n5377, C2 => 
                           MEM_IN(27), A => n5492, ZN => n5491);
   U5969 : OAI22_X1 port map( A1 => n11698, A2 => n233, B1 => n5141, B2 => 
                           n5380, ZN => n5492);
   U5970 : AOI22_X1 port map( A1 => n5381, A2 => n5142, B1 => n5382, B2 => 
                           n5143, ZN => n5490);
   U5971 : AOI22_X1 port map( A1 => n5383, A2 => n5144, B1 => n5384, B2 => 
                           n5145, ZN => n5489);
   U5972 : NAND3_X1 port map( A1 => n5493, A2 => n5494, A3 => n5495, ZN => 
                           n13060);
   U5973 : AOI221_X1 port map( B1 => n5376, B2 => n5149, C1 => n5377, C2 => 
                           MEM_IN(28), A => n5496, ZN => n5495);
   U5974 : OAI22_X1 port map( A1 => n11697, A2 => n233, B1 => n5151, B2 => 
                           n5380, ZN => n5496);
   U5975 : AOI22_X1 port map( A1 => n5381, A2 => n5152, B1 => n5382, B2 => 
                           n5153, ZN => n5494);
   U5976 : AOI22_X1 port map( A1 => n5383, A2 => n5154, B1 => n5384, B2 => 
                           n5155, ZN => n5493);
   U5977 : NAND3_X1 port map( A1 => n5497, A2 => n5498, A3 => n5499, ZN => 
                           n13059);
   U5978 : AOI221_X1 port map( B1 => n5376, B2 => n5159, C1 => n5377, C2 => 
                           MEM_IN(29), A => n5500, ZN => n5499);
   U5979 : OAI22_X1 port map( A1 => n11696, A2 => n233, B1 => n5161, B2 => 
                           n5380, ZN => n5500);
   U5980 : AOI22_X1 port map( A1 => n5381, A2 => n5162, B1 => n5382, B2 => 
                           n5163, ZN => n5498);
   U5981 : AOI22_X1 port map( A1 => n5383, A2 => n5164, B1 => n5384, B2 => 
                           n5165, ZN => n5497);
   U5982 : NAND3_X1 port map( A1 => n5501, A2 => n5502, A3 => n5503, ZN => 
                           n13058);
   U5983 : AOI221_X1 port map( B1 => n5376, B2 => n5169, C1 => n5377, C2 => 
                           MEM_IN(30), A => n5504, ZN => n5503);
   U5984 : OAI22_X1 port map( A1 => n11695, A2 => n233, B1 => n5171, B2 => 
                           n5380, ZN => n5504);
   U5985 : AOI22_X1 port map( A1 => n5381, A2 => n5172, B1 => n5382, B2 => 
                           n5173, ZN => n5502);
   U5986 : AOI22_X1 port map( A1 => n5383, A2 => n5174, B1 => n5384, B2 => 
                           n5175, ZN => n5501);
   U5987 : NAND3_X1 port map( A1 => n5505, A2 => n5506, A3 => n5507, ZN => 
                           n13057);
   U5988 : AOI221_X1 port map( B1 => n5376, B2 => n5179, C1 => n5377, C2 => 
                           MEM_IN(31), A => n5508, ZN => n5507);
   U5989 : OAI22_X1 port map( A1 => n11694, A2 => n233, B1 => n5181, B2 => 
                           n5380, ZN => n5508);
   U5990 : OAI211_X1 port map( C1 => n5513, C2 => n4787, A => n5514, B => n5515
                           , ZN => n5512);
   U5991 : AND3_X1 port map( A1 => n5198, A2 => n5516, A3 => n5369, ZN => n5513
                           );
   U5992 : INV_X1 port map( A => n5190, ZN => n5198);
   U5993 : AOI22_X1 port map( A1 => n5381, A2 => n5191, B1 => n5382, B2 => 
                           n5192, ZN => n5506);
   U5994 : AOI22_X1 port map( A1 => n5383, A2 => n5195, B1 => n5384, B2 => 
                           n5196, ZN => n5505);
   U5995 : OAI22_X1 port map( A1 => n5511, A2 => n5518, B1 => n208, B2 => n232,
                           ZN => n5514);
   U5996 : INV_X1 port map( A => n5510, ZN => n5518);
   U5997 : NOR3_X1 port map( A1 => n4841, A2 => n232, A3 => n5509, ZN => n5510)
                           ;
   U5998 : OAI22_X1 port map( A1 => n4786, A2 => n5519, B1 => n5520, B2 => 
                           n5204, ZN => n5379);
   U5999 : NOR2_X1 port map( A1 => n5509, A2 => n5511, ZN => n5520);
   U6000 : NAND2_X1 port map( A1 => n5364, A2 => n5521, ZN => n5509);
   U6001 : NOR2_X1 port map( A1 => n5211, A2 => n5214, ZN => n5364);
   U6002 : AOI221_X1 port map( B1 => n5522, B2 => n5208, C1 => n5206, C2 => 
                           n5211, A => RESET, ZN => n5519);
   U6003 : NAND2_X1 port map( A1 => n5523, A2 => n5369, ZN => n5211);
   U6004 : OR2_X1 port map( A1 => n5524, A2 => n5525, ZN => n5511);
   U6005 : NOR2_X1 port map( A1 => n5190, A2 => n5369, ZN => n5193);
   U6006 : NAND2_X1 port map( A1 => n5526, A2 => n5216, ZN => n5369);
   U6007 : NAND3_X1 port map( A1 => n5527, A2 => n5528, A3 => n5529, ZN => 
                           n13056);
   U6008 : AOI221_X1 port map( B1 => n5530, B2 => n5531, C1 => n5532, C2 => 
                           REGISTERS_36_0_port, A => n5533, ZN => n5529);
   U6009 : OAI22_X1 port map( A1 => n5534, A2 => n5535, B1 => n5536, B2 => 
                           n5537, ZN => n5533);
   U6010 : AOI22_X1 port map( A1 => n202, A2 => n4869, B1 => n167, B2 => n4871,
                           ZN => n5528);
   U6011 : AOI22_X1 port map( A1 => n203, A2 => n4873, B1 => n164, B2 => n4875,
                           ZN => n5527);
   U6012 : NAND3_X1 port map( A1 => n5538, A2 => n5539, A3 => n5540, ZN => 
                           n13055);
   U6013 : AOI221_X1 port map( B1 => n5530, B2 => n5541, C1 => n5532, C2 => 
                           REGISTERS_36_1_port, A => n5542, ZN => n5540);
   U6014 : OAI22_X1 port map( A1 => n5543, A2 => n5535, B1 => n5544, B2 => 
                           n5537, ZN => n5542);
   U6015 : AOI22_X1 port map( A1 => n202, A2 => n4882, B1 => n167, B2 => n4883,
                           ZN => n5539);
   U6016 : AOI22_X1 port map( A1 => n203, A2 => n4884, B1 => n164, B2 => n4885,
                           ZN => n5538);
   U6017 : NAND3_X1 port map( A1 => n5545, A2 => n5546, A3 => n5547, ZN => 
                           n13054);
   U6018 : AOI221_X1 port map( B1 => n5530, B2 => n5548, C1 => n5532, C2 => 
                           REGISTERS_36_2_port, A => n5549, ZN => n5547);
   U6019 : OAI22_X1 port map( A1 => n5550, A2 => n5535, B1 => n5551, B2 => 
                           n5537, ZN => n5549);
   U6020 : AOI22_X1 port map( A1 => n202, A2 => n4892, B1 => n167, B2 => n4893,
                           ZN => n5546);
   U6021 : AOI22_X1 port map( A1 => n203, A2 => n4894, B1 => n164, B2 => n4895,
                           ZN => n5545);
   U6022 : NAND3_X1 port map( A1 => n5552, A2 => n5553, A3 => n5554, ZN => 
                           n13053);
   U6023 : AOI221_X1 port map( B1 => n5530, B2 => n5555, C1 => n5532, C2 => 
                           REGISTERS_36_3_port, A => n5556, ZN => n5554);
   U6024 : OAI22_X1 port map( A1 => n5557, A2 => n5535, B1 => n5558, B2 => 
                           n5537, ZN => n5556);
   U6025 : AOI22_X1 port map( A1 => n202, A2 => n4902, B1 => n167, B2 => n4903,
                           ZN => n5553);
   U6026 : AOI22_X1 port map( A1 => n203, A2 => n4904, B1 => n164, B2 => n4905,
                           ZN => n5552);
   U6027 : NAND3_X1 port map( A1 => n5559, A2 => n5560, A3 => n5561, ZN => 
                           n13052);
   U6028 : AOI221_X1 port map( B1 => n5530, B2 => n5562, C1 => n5532, C2 => 
                           REGISTERS_36_4_port, A => n5563, ZN => n5561);
   U6029 : OAI22_X1 port map( A1 => n5564, A2 => n5535, B1 => n5565, B2 => 
                           n5537, ZN => n5563);
   U6030 : AOI22_X1 port map( A1 => n202, A2 => n4912, B1 => n167, B2 => n4913,
                           ZN => n5560);
   U6031 : AOI22_X1 port map( A1 => n203, A2 => n4914, B1 => n164, B2 => n4915,
                           ZN => n5559);
   U6032 : NAND3_X1 port map( A1 => n5566, A2 => n5567, A3 => n5568, ZN => 
                           n13051);
   U6033 : AOI221_X1 port map( B1 => n5530, B2 => n5569, C1 => n5532, C2 => 
                           REGISTERS_36_5_port, A => n5570, ZN => n5568);
   U6034 : OAI22_X1 port map( A1 => n5571, A2 => n5535, B1 => n5572, B2 => 
                           n5537, ZN => n5570);
   U6035 : AOI22_X1 port map( A1 => n202, A2 => n4922, B1 => n167, B2 => n4923,
                           ZN => n5567);
   U6036 : AOI22_X1 port map( A1 => n203, A2 => n4924, B1 => n164, B2 => n4925,
                           ZN => n5566);
   U6037 : NAND3_X1 port map( A1 => n5573, A2 => n5574, A3 => n5575, ZN => 
                           n13050);
   U6038 : AOI221_X1 port map( B1 => n5530, B2 => n5576, C1 => n5532, C2 => 
                           REGISTERS_36_6_port, A => n5577, ZN => n5575);
   U6039 : OAI22_X1 port map( A1 => n5578, A2 => n5535, B1 => n5579, B2 => 
                           n5537, ZN => n5577);
   U6040 : AOI22_X1 port map( A1 => n202, A2 => n4932, B1 => n167, B2 => n4933,
                           ZN => n5574);
   U6041 : AOI22_X1 port map( A1 => n203, A2 => n4934, B1 => n164, B2 => n4935,
                           ZN => n5573);
   U6042 : NAND3_X1 port map( A1 => n5580, A2 => n5581, A3 => n5582, ZN => 
                           n13049);
   U6043 : AOI221_X1 port map( B1 => n5530, B2 => n5583, C1 => n5532, C2 => 
                           REGISTERS_36_7_port, A => n5584, ZN => n5582);
   U6044 : OAI22_X1 port map( A1 => n5585, A2 => n5535, B1 => n5586, B2 => 
                           n5537, ZN => n5584);
   U6045 : AOI22_X1 port map( A1 => n202, A2 => n4942, B1 => n167, B2 => n4943,
                           ZN => n5581);
   U6046 : AOI22_X1 port map( A1 => n203, A2 => n4944, B1 => n164, B2 => n4945,
                           ZN => n5580);
   U6047 : NAND3_X1 port map( A1 => n5587, A2 => n5588, A3 => n5589, ZN => 
                           n13048);
   U6048 : AOI221_X1 port map( B1 => n5530, B2 => n5590, C1 => n5532, C2 => 
                           REGISTERS_36_8_port, A => n5591, ZN => n5589);
   U6049 : OAI22_X1 port map( A1 => n5592, A2 => n5535, B1 => n5593, B2 => 
                           n5537, ZN => n5591);
   U6050 : AOI22_X1 port map( A1 => n202, A2 => n4952, B1 => n167, B2 => n4953,
                           ZN => n5588);
   U6051 : AOI22_X1 port map( A1 => n203, A2 => n4954, B1 => n164, B2 => n4955,
                           ZN => n5587);
   U6052 : NAND3_X1 port map( A1 => n5594, A2 => n5595, A3 => n5596, ZN => 
                           n13047);
   U6053 : AOI221_X1 port map( B1 => n5530, B2 => n5597, C1 => n5532, C2 => 
                           REGISTERS_36_9_port, A => n5598, ZN => n5596);
   U6054 : OAI22_X1 port map( A1 => n5599, A2 => n5535, B1 => n5600, B2 => 
                           n5537, ZN => n5598);
   U6055 : AOI22_X1 port map( A1 => n202, A2 => n4962, B1 => n167, B2 => n4963,
                           ZN => n5595);
   U6056 : AOI22_X1 port map( A1 => n203, A2 => n4964, B1 => n164, B2 => n4965,
                           ZN => n5594);
   U6057 : NAND3_X1 port map( A1 => n5601, A2 => n5602, A3 => n5603, ZN => 
                           n13046);
   U6058 : AOI221_X1 port map( B1 => n5530, B2 => n5604, C1 => n5532, C2 => 
                           REGISTERS_36_10_port, A => n5605, ZN => n5603);
   U6059 : OAI22_X1 port map( A1 => n5606, A2 => n5535, B1 => n5607, B2 => 
                           n5537, ZN => n5605);
   U6060 : AOI22_X1 port map( A1 => n202, A2 => n4972, B1 => n167, B2 => n4973,
                           ZN => n5602);
   U6061 : AOI22_X1 port map( A1 => n203, A2 => n4974, B1 => n164, B2 => n4975,
                           ZN => n5601);
   U6062 : NAND3_X1 port map( A1 => n5608, A2 => n5609, A3 => n5610, ZN => 
                           n13045);
   U6063 : AOI221_X1 port map( B1 => n5530, B2 => n5611, C1 => n5532, C2 => 
                           REGISTERS_36_11_port, A => n5612, ZN => n5610);
   U6064 : OAI22_X1 port map( A1 => n5613, A2 => n5535, B1 => n5614, B2 => 
                           n5537, ZN => n5612);
   U6065 : AOI22_X1 port map( A1 => n202, A2 => n4982, B1 => n167, B2 => n4983,
                           ZN => n5609);
   U6066 : AOI22_X1 port map( A1 => n203, A2 => n4984, B1 => n164, B2 => n4985,
                           ZN => n5608);
   U6067 : NAND3_X1 port map( A1 => n5615, A2 => n5616, A3 => n5617, ZN => 
                           n13044);
   U6068 : AOI221_X1 port map( B1 => n5530, B2 => n5618, C1 => n5532, C2 => 
                           REGISTERS_36_12_port, A => n5619, ZN => n5617);
   U6069 : OAI22_X1 port map( A1 => n5620, A2 => n5535, B1 => n5621, B2 => 
                           n5537, ZN => n5619);
   U6070 : AOI22_X1 port map( A1 => n202, A2 => n4992, B1 => n167, B2 => n4993,
                           ZN => n5616);
   U6071 : AOI22_X1 port map( A1 => n203, A2 => n4994, B1 => n164, B2 => n4995,
                           ZN => n5615);
   U6072 : NAND3_X1 port map( A1 => n5622, A2 => n5623, A3 => n5624, ZN => 
                           n13043);
   U6073 : AOI221_X1 port map( B1 => n5530, B2 => n5625, C1 => n5532, C2 => 
                           REGISTERS_36_13_port, A => n5626, ZN => n5624);
   U6074 : OAI22_X1 port map( A1 => n5627, A2 => n5535, B1 => n5628, B2 => 
                           n5537, ZN => n5626);
   U6075 : AOI22_X1 port map( A1 => n202, A2 => n5002, B1 => n167, B2 => n5003,
                           ZN => n5623);
   U6076 : AOI22_X1 port map( A1 => n203, A2 => n5004, B1 => n164, B2 => n5005,
                           ZN => n5622);
   U6077 : NAND3_X1 port map( A1 => n5629, A2 => n5630, A3 => n5631, ZN => 
                           n13042);
   U6078 : AOI221_X1 port map( B1 => n5530, B2 => n5632, C1 => n5532, C2 => 
                           REGISTERS_36_14_port, A => n5633, ZN => n5631);
   U6079 : OAI22_X1 port map( A1 => n5634, A2 => n5535, B1 => n5635, B2 => 
                           n5537, ZN => n5633);
   U6080 : AOI22_X1 port map( A1 => n202, A2 => n5012, B1 => n167, B2 => n5013,
                           ZN => n5630);
   U6081 : AOI22_X1 port map( A1 => n203, A2 => n5014, B1 => n164, B2 => n5015,
                           ZN => n5629);
   U6082 : NAND3_X1 port map( A1 => n5636, A2 => n5637, A3 => n5638, ZN => 
                           n13041);
   U6083 : AOI221_X1 port map( B1 => n5530, B2 => n5639, C1 => n5532, C2 => 
                           REGISTERS_36_15_port, A => n5640, ZN => n5638);
   U6084 : OAI22_X1 port map( A1 => n5641, A2 => n5535, B1 => n5642, B2 => 
                           n5537, ZN => n5640);
   U6085 : AOI22_X1 port map( A1 => n202, A2 => n5022, B1 => n167, B2 => n5023,
                           ZN => n5637);
   U6086 : AOI22_X1 port map( A1 => n203, A2 => n5024, B1 => n164, B2 => n5025,
                           ZN => n5636);
   U6087 : NAND3_X1 port map( A1 => n5643, A2 => n5644, A3 => n5645, ZN => 
                           n13040);
   U6088 : AOI221_X1 port map( B1 => n5530, B2 => n5646, C1 => n5532, C2 => 
                           REGISTERS_36_16_port, A => n5647, ZN => n5645);
   U6089 : OAI22_X1 port map( A1 => n5648, A2 => n5535, B1 => n5649, B2 => 
                           n5537, ZN => n5647);
   U6090 : AOI22_X1 port map( A1 => n202, A2 => n5032, B1 => n167, B2 => n5033,
                           ZN => n5644);
   U6091 : AOI22_X1 port map( A1 => n203, A2 => n5034, B1 => n164, B2 => n5035,
                           ZN => n5643);
   U6092 : NAND3_X1 port map( A1 => n5650, A2 => n5651, A3 => n5652, ZN => 
                           n13039);
   U6093 : AOI221_X1 port map( B1 => n5530, B2 => n5653, C1 => n5532, C2 => 
                           REGISTERS_36_17_port, A => n5654, ZN => n5652);
   U6094 : OAI22_X1 port map( A1 => n5655, A2 => n5535, B1 => n5656, B2 => 
                           n5537, ZN => n5654);
   U6095 : AOI22_X1 port map( A1 => n202, A2 => n5042, B1 => n167, B2 => n5043,
                           ZN => n5651);
   U6096 : AOI22_X1 port map( A1 => n203, A2 => n5044, B1 => n164, B2 => n5045,
                           ZN => n5650);
   U6097 : NAND3_X1 port map( A1 => n5657, A2 => n5658, A3 => n5659, ZN => 
                           n13038);
   U6098 : AOI221_X1 port map( B1 => n5530, B2 => n5660, C1 => n5532, C2 => 
                           REGISTERS_36_18_port, A => n5661, ZN => n5659);
   U6099 : OAI22_X1 port map( A1 => n5662, A2 => n5535, B1 => n5663, B2 => 
                           n5537, ZN => n5661);
   U6100 : AOI22_X1 port map( A1 => n202, A2 => n5052, B1 => n167, B2 => n5053,
                           ZN => n5658);
   U6101 : AOI22_X1 port map( A1 => n203, A2 => n5054, B1 => n164, B2 => n5055,
                           ZN => n5657);
   U6102 : NAND3_X1 port map( A1 => n5664, A2 => n5665, A3 => n5666, ZN => 
                           n13037);
   U6103 : AOI221_X1 port map( B1 => n5530, B2 => n5667, C1 => n5532, C2 => 
                           REGISTERS_36_19_port, A => n5668, ZN => n5666);
   U6104 : OAI22_X1 port map( A1 => n5669, A2 => n5535, B1 => n5670, B2 => 
                           n5537, ZN => n5668);
   U6105 : AOI22_X1 port map( A1 => n202, A2 => n5062, B1 => n167, B2 => n5063,
                           ZN => n5665);
   U6106 : AOI22_X1 port map( A1 => n203, A2 => n5064, B1 => n164, B2 => n5065,
                           ZN => n5664);
   U6107 : NAND3_X1 port map( A1 => n5671, A2 => n5672, A3 => n5673, ZN => 
                           n13036);
   U6108 : AOI221_X1 port map( B1 => n5530, B2 => n5674, C1 => n5532, C2 => 
                           REGISTERS_36_20_port, A => n5675, ZN => n5673);
   U6109 : OAI22_X1 port map( A1 => n5676, A2 => n5535, B1 => n5677, B2 => 
                           n5537, ZN => n5675);
   U6110 : AOI22_X1 port map( A1 => n202, A2 => n5072, B1 => n167, B2 => n5073,
                           ZN => n5672);
   U6111 : AOI22_X1 port map( A1 => n203, A2 => n5074, B1 => n164, B2 => n5075,
                           ZN => n5671);
   U6112 : NAND3_X1 port map( A1 => n5678, A2 => n5679, A3 => n5680, ZN => 
                           n13035);
   U6113 : AOI221_X1 port map( B1 => n5530, B2 => n5681, C1 => n5532, C2 => 
                           REGISTERS_36_21_port, A => n5682, ZN => n5680);
   U6114 : OAI22_X1 port map( A1 => n5683, A2 => n5535, B1 => n5684, B2 => 
                           n5537, ZN => n5682);
   U6115 : AOI22_X1 port map( A1 => n202, A2 => n5082, B1 => n167, B2 => n5083,
                           ZN => n5679);
   U6116 : AOI22_X1 port map( A1 => n203, A2 => n5084, B1 => n164, B2 => n5085,
                           ZN => n5678);
   U6117 : NAND3_X1 port map( A1 => n5685, A2 => n5686, A3 => n5687, ZN => 
                           n13034);
   U6118 : AOI221_X1 port map( B1 => n5530, B2 => n5688, C1 => n5532, C2 => 
                           REGISTERS_36_22_port, A => n5689, ZN => n5687);
   U6119 : OAI22_X1 port map( A1 => n5690, A2 => n5535, B1 => n5691, B2 => 
                           n5537, ZN => n5689);
   U6120 : AOI22_X1 port map( A1 => n202, A2 => n5092, B1 => n167, B2 => n5093,
                           ZN => n5686);
   U6121 : AOI22_X1 port map( A1 => n203, A2 => n5094, B1 => n164, B2 => n5095,
                           ZN => n5685);
   U6122 : NAND3_X1 port map( A1 => n5692, A2 => n5693, A3 => n5694, ZN => 
                           n13033);
   U6123 : AOI221_X1 port map( B1 => n5530, B2 => n5695, C1 => n5532, C2 => 
                           REGISTERS_36_23_port, A => n5696, ZN => n5694);
   U6124 : OAI22_X1 port map( A1 => n5697, A2 => n5535, B1 => n5698, B2 => 
                           n5537, ZN => n5696);
   U6125 : AOI22_X1 port map( A1 => n202, A2 => n5102, B1 => n167, B2 => n5103,
                           ZN => n5693);
   U6126 : AOI22_X1 port map( A1 => n203, A2 => n5104, B1 => n164, B2 => n5105,
                           ZN => n5692);
   U6127 : NAND3_X1 port map( A1 => n5699, A2 => n5700, A3 => n5701, ZN => 
                           n13032);
   U6128 : AOI221_X1 port map( B1 => n5530, B2 => n5702, C1 => n5532, C2 => 
                           REGISTERS_36_24_port, A => n5703, ZN => n5701);
   U6129 : OAI22_X1 port map( A1 => n5704, A2 => n5535, B1 => n5705, B2 => 
                           n5537, ZN => n5703);
   U6130 : AOI22_X1 port map( A1 => n202, A2 => n5112, B1 => n167, B2 => n5113,
                           ZN => n5700);
   U6131 : AOI22_X1 port map( A1 => n203, A2 => n5114, B1 => n164, B2 => n5115,
                           ZN => n5699);
   U6132 : NAND3_X1 port map( A1 => n5706, A2 => n5707, A3 => n5708, ZN => 
                           n13031);
   U6133 : AOI221_X1 port map( B1 => n5530, B2 => n5709, C1 => n5532, C2 => 
                           REGISTERS_36_25_port, A => n5710, ZN => n5708);
   U6134 : OAI22_X1 port map( A1 => n5711, A2 => n5535, B1 => n5712, B2 => 
                           n5537, ZN => n5710);
   U6135 : AOI22_X1 port map( A1 => n202, A2 => n5122, B1 => n167, B2 => n5123,
                           ZN => n5707);
   U6136 : AOI22_X1 port map( A1 => n203, A2 => n5124, B1 => n164, B2 => n5125,
                           ZN => n5706);
   U6137 : NAND3_X1 port map( A1 => n5713, A2 => n5714, A3 => n5715, ZN => 
                           n13030);
   U6138 : AOI221_X1 port map( B1 => n5530, B2 => n5716, C1 => n5532, C2 => 
                           REGISTERS_36_26_port, A => n5717, ZN => n5715);
   U6139 : OAI22_X1 port map( A1 => n5718, A2 => n5535, B1 => n5719, B2 => 
                           n5537, ZN => n5717);
   U6140 : AOI22_X1 port map( A1 => n202, A2 => n5132, B1 => n167, B2 => n5133,
                           ZN => n5714);
   U6141 : AOI22_X1 port map( A1 => n203, A2 => n5134, B1 => n164, B2 => n5135,
                           ZN => n5713);
   U6142 : NAND3_X1 port map( A1 => n5720, A2 => n5721, A3 => n5722, ZN => 
                           n13029);
   U6143 : AOI221_X1 port map( B1 => n5530, B2 => n5723, C1 => n5532, C2 => 
                           REGISTERS_36_27_port, A => n5724, ZN => n5722);
   U6144 : OAI22_X1 port map( A1 => n5725, A2 => n5535, B1 => n5726, B2 => 
                           n5537, ZN => n5724);
   U6145 : AOI22_X1 port map( A1 => n202, A2 => n5142, B1 => n167, B2 => n5143,
                           ZN => n5721);
   U6146 : AOI22_X1 port map( A1 => n203, A2 => n5144, B1 => n164, B2 => n5145,
                           ZN => n5720);
   U6147 : NAND3_X1 port map( A1 => n5727, A2 => n5728, A3 => n5729, ZN => 
                           n13028);
   U6148 : AOI221_X1 port map( B1 => n5530, B2 => n5730, C1 => n5532, C2 => 
                           REGISTERS_36_28_port, A => n5731, ZN => n5729);
   U6149 : OAI22_X1 port map( A1 => n5732, A2 => n5535, B1 => n5733, B2 => 
                           n5537, ZN => n5731);
   U6150 : AOI22_X1 port map( A1 => n202, A2 => n5152, B1 => n167, B2 => n5153,
                           ZN => n5728);
   U6151 : AOI22_X1 port map( A1 => n203, A2 => n5154, B1 => n164, B2 => n5155,
                           ZN => n5727);
   U6152 : NAND3_X1 port map( A1 => n5734, A2 => n5735, A3 => n5736, ZN => 
                           n13027);
   U6153 : AOI221_X1 port map( B1 => n5530, B2 => n5737, C1 => n5532, C2 => 
                           REGISTERS_36_29_port, A => n5738, ZN => n5736);
   U6154 : OAI22_X1 port map( A1 => n5739, A2 => n5535, B1 => n5740, B2 => 
                           n5537, ZN => n5738);
   U6155 : AOI22_X1 port map( A1 => n202, A2 => n5162, B1 => n167, B2 => n5163,
                           ZN => n5735);
   U6156 : AOI22_X1 port map( A1 => n203, A2 => n5164, B1 => n164, B2 => n5165,
                           ZN => n5734);
   U6157 : NAND3_X1 port map( A1 => n5741, A2 => n5742, A3 => n5743, ZN => 
                           n13026);
   U6158 : AOI221_X1 port map( B1 => n5530, B2 => n5744, C1 => n5532, C2 => 
                           REGISTERS_36_30_port, A => n5745, ZN => n5743);
   U6159 : OAI22_X1 port map( A1 => n5746, A2 => n5535, B1 => n5747, B2 => 
                           n5537, ZN => n5745);
   U6160 : AOI22_X1 port map( A1 => n202, A2 => n5172, B1 => n167, B2 => n5173,
                           ZN => n5742);
   U6161 : AOI22_X1 port map( A1 => n203, A2 => n5174, B1 => n164, B2 => n5175,
                           ZN => n5741);
   U6162 : NAND3_X1 port map( A1 => n5748, A2 => n5749, A3 => n5750, ZN => 
                           n13025);
   U6163 : AOI221_X1 port map( B1 => n5530, B2 => n5751, C1 => n5532, C2 => 
                           REGISTERS_36_31_port, A => n5752, ZN => n5750);
   U6164 : OAI22_X1 port map( A1 => n5753, A2 => n5535, B1 => n5754, B2 => 
                           n5537, ZN => n5752);
   U6165 : AOI21_X1 port map( B1 => n5206, B2 => n5190, A => n5758, ZN => n5757
                           );
   U6166 : NAND2_X1 port map( A1 => n5206, A2 => n5759, ZN => n5190);
   U6167 : AOI22_X1 port map( A1 => n202, A2 => n5191, B1 => n167, B2 => n5192,
                           ZN => n5749);
   U6168 : AOI22_X1 port map( A1 => n203, A2 => n5195, B1 => n164, B2 => n5196,
                           ZN => n5748);
   U6169 : AOI22_X1 port map( A1 => n5764, A2 => n5760, B1 => n4841, B2 => 
                           n5762, ZN => n5758);
   U6170 : NOR3_X1 port map( A1 => n4841, A2 => n5532, A3 => n5763, ZN => n5760
                           );
   U6171 : OAI22_X1 port map( A1 => n4786, A2 => n5765, B1 => n5766, B2 => 
                           n5204, ZN => n5762);
   U6172 : NOR2_X1 port map( A1 => n5763, A2 => n5761, ZN => n5766);
   U6173 : NAND2_X1 port map( A1 => n5767, A2 => n5523, ZN => n5763);
   U6174 : NOR3_X1 port map( A1 => n5768, A2 => RESET, A3 => n5769, ZN => n5765
                           );
   U6175 : OAI22_X1 port map( A1 => n5770, A2 => n5771, B1 => n5523, B2 => 
                           n4787, ZN => n5768);
   U6176 : AND3_X1 port map( A1 => n5516, A2 => n5772, A3 => n5759, ZN => n5523
                           );
   U6177 : INV_X1 port map( A => n5761, ZN => n5764);
   U6178 : NAND2_X1 port map( A1 => n5773, A2 => n5774, ZN => n5761);
   U6179 : INV_X1 port map( A => n5194, ZN => n5367);
   U6180 : NOR2_X1 port map( A1 => n5759, A2 => n4787, ZN => n5194);
   U6181 : NAND2_X1 port map( A1 => n5775, A2 => n5216, ZN => n5759);
   U6182 : NAND3_X1 port map( A1 => n5776, A2 => n5777, A3 => n5778, ZN => 
                           n13024);
   U6183 : AOI221_X1 port map( B1 => n5779, B2 => n4863, C1 => n5780, C2 => 
                           MEM_IN(0), A => n5781, ZN => n5778);
   U6184 : OAI22_X1 port map( A1 => n11661, A2 => n235, B1 => n4867, B2 => 
                           n5783, ZN => n5781);
   U6185 : AOI22_X1 port map( A1 => n5784, A2 => n4869, B1 => n5785, B2 => 
                           n4871, ZN => n5777);
   U6186 : AOI22_X1 port map( A1 => n5786, A2 => n4873, B1 => n5787, B2 => 
                           n4875, ZN => n5776);
   U6187 : NAND3_X1 port map( A1 => n5788, A2 => n5789, A3 => n5790, ZN => 
                           n13023);
   U6188 : AOI221_X1 port map( B1 => n5779, B2 => n4879, C1 => n5780, C2 => 
                           MEM_IN(1), A => n5791, ZN => n5790);
   U6189 : OAI22_X1 port map( A1 => n11660, A2 => n235, B1 => n4881, B2 => 
                           n5783, ZN => n5791);
   U6190 : AOI22_X1 port map( A1 => n5784, A2 => n4882, B1 => n5785, B2 => 
                           n4883, ZN => n5789);
   U6191 : AOI22_X1 port map( A1 => n5786, A2 => n4884, B1 => n5787, B2 => 
                           n4885, ZN => n5788);
   U6192 : NAND3_X1 port map( A1 => n5792, A2 => n5793, A3 => n5794, ZN => 
                           n13022);
   U6193 : AOI221_X1 port map( B1 => n5779, B2 => n4889, C1 => n5780, C2 => 
                           MEM_IN(2), A => n5795, ZN => n5794);
   U6194 : OAI22_X1 port map( A1 => n11659, A2 => n235, B1 => n4891, B2 => 
                           n5783, ZN => n5795);
   U6195 : AOI22_X1 port map( A1 => n5784, A2 => n4892, B1 => n5785, B2 => 
                           n4893, ZN => n5793);
   U6196 : AOI22_X1 port map( A1 => n5786, A2 => n4894, B1 => n5787, B2 => 
                           n4895, ZN => n5792);
   U6197 : NAND3_X1 port map( A1 => n5796, A2 => n5797, A3 => n5798, ZN => 
                           n13021);
   U6198 : AOI221_X1 port map( B1 => n5779, B2 => n4899, C1 => n5780, C2 => 
                           MEM_IN(3), A => n5799, ZN => n5798);
   U6199 : OAI22_X1 port map( A1 => n11658, A2 => n235, B1 => n4901, B2 => 
                           n5783, ZN => n5799);
   U6200 : AOI22_X1 port map( A1 => n5784, A2 => n4902, B1 => n5785, B2 => 
                           n4903, ZN => n5797);
   U6201 : AOI22_X1 port map( A1 => n5786, A2 => n4904, B1 => n5787, B2 => 
                           n4905, ZN => n5796);
   U6202 : NAND3_X1 port map( A1 => n5800, A2 => n5801, A3 => n5802, ZN => 
                           n13020);
   U6203 : AOI221_X1 port map( B1 => n5779, B2 => n4909, C1 => n5780, C2 => 
                           MEM_IN(4), A => n5803, ZN => n5802);
   U6204 : OAI22_X1 port map( A1 => n11657, A2 => n235, B1 => n4911, B2 => 
                           n5783, ZN => n5803);
   U6205 : AOI22_X1 port map( A1 => n5784, A2 => n4912, B1 => n5785, B2 => 
                           n4913, ZN => n5801);
   U6206 : AOI22_X1 port map( A1 => n5786, A2 => n4914, B1 => n5787, B2 => 
                           n4915, ZN => n5800);
   U6207 : NAND3_X1 port map( A1 => n5804, A2 => n5805, A3 => n5806, ZN => 
                           n13019);
   U6208 : AOI221_X1 port map( B1 => n5779, B2 => n4919, C1 => n5780, C2 => 
                           MEM_IN(5), A => n5807, ZN => n5806);
   U6209 : OAI22_X1 port map( A1 => n11656, A2 => n235, B1 => n4921, B2 => 
                           n5783, ZN => n5807);
   U6210 : AOI22_X1 port map( A1 => n5784, A2 => n4922, B1 => n5785, B2 => 
                           n4923, ZN => n5805);
   U6211 : AOI22_X1 port map( A1 => n5786, A2 => n4924, B1 => n5787, B2 => 
                           n4925, ZN => n5804);
   U6212 : NAND3_X1 port map( A1 => n5808, A2 => n5809, A3 => n5810, ZN => 
                           n13018);
   U6213 : AOI221_X1 port map( B1 => n5779, B2 => n4929, C1 => n5780, C2 => 
                           MEM_IN(6), A => n5811, ZN => n5810);
   U6214 : OAI22_X1 port map( A1 => n11655, A2 => n235, B1 => n4931, B2 => 
                           n5783, ZN => n5811);
   U6215 : AOI22_X1 port map( A1 => n5784, A2 => n4932, B1 => n5785, B2 => 
                           n4933, ZN => n5809);
   U6216 : AOI22_X1 port map( A1 => n5786, A2 => n4934, B1 => n5787, B2 => 
                           n4935, ZN => n5808);
   U6217 : NAND3_X1 port map( A1 => n5812, A2 => n5813, A3 => n5814, ZN => 
                           n13017);
   U6218 : AOI221_X1 port map( B1 => n5779, B2 => n4939, C1 => n5780, C2 => 
                           MEM_IN(7), A => n5815, ZN => n5814);
   U6219 : OAI22_X1 port map( A1 => n11654, A2 => n235, B1 => n4941, B2 => 
                           n5783, ZN => n5815);
   U6220 : AOI22_X1 port map( A1 => n5784, A2 => n4942, B1 => n5785, B2 => 
                           n4943, ZN => n5813);
   U6221 : AOI22_X1 port map( A1 => n5786, A2 => n4944, B1 => n5787, B2 => 
                           n4945, ZN => n5812);
   U6222 : NAND3_X1 port map( A1 => n5816, A2 => n5817, A3 => n5818, ZN => 
                           n13016);
   U6223 : AOI221_X1 port map( B1 => n5779, B2 => n4949, C1 => n5780, C2 => 
                           MEM_IN(8), A => n5819, ZN => n5818);
   U6224 : OAI22_X1 port map( A1 => n11653, A2 => n235, B1 => n4951, B2 => 
                           n5783, ZN => n5819);
   U6225 : AOI22_X1 port map( A1 => n5784, A2 => n4952, B1 => n5785, B2 => 
                           n4953, ZN => n5817);
   U6226 : AOI22_X1 port map( A1 => n5786, A2 => n4954, B1 => n5787, B2 => 
                           n4955, ZN => n5816);
   U6227 : NAND3_X1 port map( A1 => n5820, A2 => n5821, A3 => n5822, ZN => 
                           n13015);
   U6228 : AOI221_X1 port map( B1 => n5779, B2 => n4959, C1 => n5780, C2 => 
                           MEM_IN(9), A => n5823, ZN => n5822);
   U6229 : OAI22_X1 port map( A1 => n11652, A2 => n235, B1 => n4961, B2 => 
                           n5783, ZN => n5823);
   U6230 : AOI22_X1 port map( A1 => n5784, A2 => n4962, B1 => n5785, B2 => 
                           n4963, ZN => n5821);
   U6231 : AOI22_X1 port map( A1 => n5786, A2 => n4964, B1 => n5787, B2 => 
                           n4965, ZN => n5820);
   U6232 : NAND3_X1 port map( A1 => n5824, A2 => n5825, A3 => n5826, ZN => 
                           n13014);
   U6233 : AOI221_X1 port map( B1 => n5779, B2 => n4969, C1 => n5780, C2 => 
                           MEM_IN(10), A => n5827, ZN => n5826);
   U6234 : OAI22_X1 port map( A1 => n11651, A2 => n235, B1 => n4971, B2 => 
                           n5783, ZN => n5827);
   U6235 : AOI22_X1 port map( A1 => n5784, A2 => n4972, B1 => n5785, B2 => 
                           n4973, ZN => n5825);
   U6236 : AOI22_X1 port map( A1 => n5786, A2 => n4974, B1 => n5787, B2 => 
                           n4975, ZN => n5824);
   U6237 : NAND3_X1 port map( A1 => n5828, A2 => n5829, A3 => n5830, ZN => 
                           n13013);
   U6238 : AOI221_X1 port map( B1 => n5779, B2 => n4979, C1 => n5780, C2 => 
                           MEM_IN(11), A => n5831, ZN => n5830);
   U6239 : OAI22_X1 port map( A1 => n11650, A2 => n235, B1 => n4981, B2 => 
                           n5783, ZN => n5831);
   U6240 : AOI22_X1 port map( A1 => n5784, A2 => n4982, B1 => n5785, B2 => 
                           n4983, ZN => n5829);
   U6241 : AOI22_X1 port map( A1 => n5786, A2 => n4984, B1 => n5787, B2 => 
                           n4985, ZN => n5828);
   U6242 : NAND3_X1 port map( A1 => n5832, A2 => n5833, A3 => n5834, ZN => 
                           n13012);
   U6243 : AOI221_X1 port map( B1 => n5779, B2 => n4989, C1 => n5780, C2 => 
                           MEM_IN(12), A => n5835, ZN => n5834);
   U6244 : OAI22_X1 port map( A1 => n11649, A2 => n235, B1 => n4991, B2 => 
                           n5783, ZN => n5835);
   U6245 : AOI22_X1 port map( A1 => n5784, A2 => n4992, B1 => n5785, B2 => 
                           n4993, ZN => n5833);
   U6246 : AOI22_X1 port map( A1 => n5786, A2 => n4994, B1 => n5787, B2 => 
                           n4995, ZN => n5832);
   U6247 : NAND3_X1 port map( A1 => n5836, A2 => n5837, A3 => n5838, ZN => 
                           n13011);
   U6248 : AOI221_X1 port map( B1 => n5779, B2 => n4999, C1 => n5780, C2 => 
                           MEM_IN(13), A => n5839, ZN => n5838);
   U6249 : OAI22_X1 port map( A1 => n11648, A2 => n235, B1 => n5001, B2 => 
                           n5783, ZN => n5839);
   U6250 : AOI22_X1 port map( A1 => n5784, A2 => n5002, B1 => n5785, B2 => 
                           n5003, ZN => n5837);
   U6251 : AOI22_X1 port map( A1 => n5786, A2 => n5004, B1 => n5787, B2 => 
                           n5005, ZN => n5836);
   U6252 : NAND3_X1 port map( A1 => n5840, A2 => n5841, A3 => n5842, ZN => 
                           n13010);
   U6253 : AOI221_X1 port map( B1 => n5779, B2 => n5009, C1 => n5780, C2 => 
                           MEM_IN(14), A => n5843, ZN => n5842);
   U6254 : OAI22_X1 port map( A1 => n11647, A2 => n235, B1 => n5011, B2 => 
                           n5783, ZN => n5843);
   U6255 : AOI22_X1 port map( A1 => n5784, A2 => n5012, B1 => n5785, B2 => 
                           n5013, ZN => n5841);
   U6256 : AOI22_X1 port map( A1 => n5786, A2 => n5014, B1 => n5787, B2 => 
                           n5015, ZN => n5840);
   U6257 : NAND3_X1 port map( A1 => n5844, A2 => n5845, A3 => n5846, ZN => 
                           n13009);
   U6258 : AOI221_X1 port map( B1 => n5779, B2 => n5019, C1 => n5780, C2 => 
                           MEM_IN(15), A => n5847, ZN => n5846);
   U6259 : OAI22_X1 port map( A1 => n11646, A2 => n235, B1 => n5021, B2 => 
                           n5783, ZN => n5847);
   U6260 : AOI22_X1 port map( A1 => n5784, A2 => n5022, B1 => n5785, B2 => 
                           n5023, ZN => n5845);
   U6261 : AOI22_X1 port map( A1 => n5786, A2 => n5024, B1 => n5787, B2 => 
                           n5025, ZN => n5844);
   U6262 : NAND3_X1 port map( A1 => n5848, A2 => n5849, A3 => n5850, ZN => 
                           n13008);
   U6263 : AOI221_X1 port map( B1 => n5779, B2 => n5029, C1 => n5780, C2 => 
                           MEM_IN(16), A => n5851, ZN => n5850);
   U6264 : OAI22_X1 port map( A1 => n11645, A2 => n235, B1 => n5031, B2 => 
                           n5783, ZN => n5851);
   U6265 : AOI22_X1 port map( A1 => n5784, A2 => n5032, B1 => n5785, B2 => 
                           n5033, ZN => n5849);
   U6266 : AOI22_X1 port map( A1 => n5786, A2 => n5034, B1 => n5787, B2 => 
                           n5035, ZN => n5848);
   U6267 : NAND3_X1 port map( A1 => n5852, A2 => n5853, A3 => n5854, ZN => 
                           n13007);
   U6268 : AOI221_X1 port map( B1 => n5779, B2 => n5039, C1 => n5780, C2 => 
                           MEM_IN(17), A => n5855, ZN => n5854);
   U6269 : OAI22_X1 port map( A1 => n11644, A2 => n235, B1 => n5041, B2 => 
                           n5783, ZN => n5855);
   U6270 : AOI22_X1 port map( A1 => n5784, A2 => n5042, B1 => n5785, B2 => 
                           n5043, ZN => n5853);
   U6271 : AOI22_X1 port map( A1 => n5786, A2 => n5044, B1 => n5787, B2 => 
                           n5045, ZN => n5852);
   U6272 : NAND3_X1 port map( A1 => n5856, A2 => n5857, A3 => n5858, ZN => 
                           n13006);
   U6273 : AOI221_X1 port map( B1 => n5779, B2 => n5049, C1 => n5780, C2 => 
                           MEM_IN(18), A => n5859, ZN => n5858);
   U6274 : OAI22_X1 port map( A1 => n11643, A2 => n235, B1 => n5051, B2 => 
                           n5783, ZN => n5859);
   U6275 : AOI22_X1 port map( A1 => n5784, A2 => n5052, B1 => n5785, B2 => 
                           n5053, ZN => n5857);
   U6276 : AOI22_X1 port map( A1 => n5786, A2 => n5054, B1 => n5787, B2 => 
                           n5055, ZN => n5856);
   U6277 : NAND3_X1 port map( A1 => n5860, A2 => n5861, A3 => n5862, ZN => 
                           n13005);
   U6278 : AOI221_X1 port map( B1 => n5779, B2 => n5059, C1 => n5780, C2 => 
                           MEM_IN(19), A => n5863, ZN => n5862);
   U6279 : OAI22_X1 port map( A1 => n11642, A2 => n235, B1 => n5061, B2 => 
                           n5783, ZN => n5863);
   U6280 : AOI22_X1 port map( A1 => n5784, A2 => n5062, B1 => n5785, B2 => 
                           n5063, ZN => n5861);
   U6281 : AOI22_X1 port map( A1 => n5786, A2 => n5064, B1 => n5787, B2 => 
                           n5065, ZN => n5860);
   U6282 : NAND3_X1 port map( A1 => n5864, A2 => n5865, A3 => n5866, ZN => 
                           n13004);
   U6283 : AOI221_X1 port map( B1 => n5779, B2 => n5069, C1 => n5780, C2 => 
                           MEM_IN(20), A => n5867, ZN => n5866);
   U6284 : OAI22_X1 port map( A1 => n11641, A2 => n235, B1 => n5071, B2 => 
                           n5783, ZN => n5867);
   U6285 : AOI22_X1 port map( A1 => n5784, A2 => n5072, B1 => n5785, B2 => 
                           n5073, ZN => n5865);
   U6286 : AOI22_X1 port map( A1 => n5786, A2 => n5074, B1 => n5787, B2 => 
                           n5075, ZN => n5864);
   U6287 : NAND3_X1 port map( A1 => n5868, A2 => n5869, A3 => n5870, ZN => 
                           n13003);
   U6288 : AOI221_X1 port map( B1 => n5779, B2 => n5079, C1 => n5780, C2 => 
                           MEM_IN(21), A => n5871, ZN => n5870);
   U6289 : OAI22_X1 port map( A1 => n11640, A2 => n235, B1 => n5081, B2 => 
                           n5783, ZN => n5871);
   U6290 : AOI22_X1 port map( A1 => n5784, A2 => n5082, B1 => n5785, B2 => 
                           n5083, ZN => n5869);
   U6291 : AOI22_X1 port map( A1 => n5786, A2 => n5084, B1 => n5787, B2 => 
                           n5085, ZN => n5868);
   U6292 : NAND3_X1 port map( A1 => n5872, A2 => n5873, A3 => n5874, ZN => 
                           n13002);
   U6293 : AOI221_X1 port map( B1 => n5779, B2 => n5089, C1 => n5780, C2 => 
                           MEM_IN(22), A => n5875, ZN => n5874);
   U6294 : OAI22_X1 port map( A1 => n11639, A2 => n235, B1 => n5091, B2 => 
                           n5783, ZN => n5875);
   U6295 : AOI22_X1 port map( A1 => n5784, A2 => n5092, B1 => n5785, B2 => 
                           n5093, ZN => n5873);
   U6296 : AOI22_X1 port map( A1 => n5786, A2 => n5094, B1 => n5787, B2 => 
                           n5095, ZN => n5872);
   U6297 : NAND3_X1 port map( A1 => n5876, A2 => n5877, A3 => n5878, ZN => 
                           n13001);
   U6298 : AOI221_X1 port map( B1 => n5779, B2 => n5099, C1 => n5780, C2 => 
                           MEM_IN(23), A => n5879, ZN => n5878);
   U6299 : OAI22_X1 port map( A1 => n11638, A2 => n235, B1 => n5101, B2 => 
                           n5783, ZN => n5879);
   U6300 : AOI22_X1 port map( A1 => n5784, A2 => n5102, B1 => n5785, B2 => 
                           n5103, ZN => n5877);
   U6301 : AOI22_X1 port map( A1 => n5786, A2 => n5104, B1 => n5787, B2 => 
                           n5105, ZN => n5876);
   U6302 : NAND3_X1 port map( A1 => n5880, A2 => n5881, A3 => n5882, ZN => 
                           n13000);
   U6303 : AOI221_X1 port map( B1 => n5779, B2 => n5109, C1 => n5780, C2 => 
                           MEM_IN(24), A => n5883, ZN => n5882);
   U6304 : OAI22_X1 port map( A1 => n11637, A2 => n235, B1 => n5111, B2 => 
                           n5783, ZN => n5883);
   U6305 : AOI22_X1 port map( A1 => n5784, A2 => n5112, B1 => n5785, B2 => 
                           n5113, ZN => n5881);
   U6306 : AOI22_X1 port map( A1 => n5786, A2 => n5114, B1 => n5787, B2 => 
                           n5115, ZN => n5880);
   U6307 : NAND3_X1 port map( A1 => n5884, A2 => n5885, A3 => n5886, ZN => 
                           n12999);
   U6308 : AOI221_X1 port map( B1 => n5779, B2 => n5119, C1 => n5780, C2 => 
                           MEM_IN(25), A => n5887, ZN => n5886);
   U6309 : OAI22_X1 port map( A1 => n11636, A2 => n235, B1 => n5121, B2 => 
                           n5783, ZN => n5887);
   U6310 : AOI22_X1 port map( A1 => n5784, A2 => n5122, B1 => n5785, B2 => 
                           n5123, ZN => n5885);
   U6311 : AOI22_X1 port map( A1 => n5786, A2 => n5124, B1 => n5787, B2 => 
                           n5125, ZN => n5884);
   U6312 : NAND3_X1 port map( A1 => n5888, A2 => n5889, A3 => n5890, ZN => 
                           n12998);
   U6313 : AOI221_X1 port map( B1 => n5779, B2 => n5129, C1 => n5780, C2 => 
                           MEM_IN(26), A => n5891, ZN => n5890);
   U6314 : OAI22_X1 port map( A1 => n11635, A2 => n235, B1 => n5131, B2 => 
                           n5783, ZN => n5891);
   U6315 : AOI22_X1 port map( A1 => n5784, A2 => n5132, B1 => n5785, B2 => 
                           n5133, ZN => n5889);
   U6316 : AOI22_X1 port map( A1 => n5786, A2 => n5134, B1 => n5787, B2 => 
                           n5135, ZN => n5888);
   U6317 : NAND3_X1 port map( A1 => n5892, A2 => n5893, A3 => n5894, ZN => 
                           n12997);
   U6318 : AOI221_X1 port map( B1 => n5779, B2 => n5139, C1 => n5780, C2 => 
                           MEM_IN(27), A => n5895, ZN => n5894);
   U6319 : OAI22_X1 port map( A1 => n11634, A2 => n235, B1 => n5141, B2 => 
                           n5783, ZN => n5895);
   U6320 : AOI22_X1 port map( A1 => n5784, A2 => n5142, B1 => n5785, B2 => 
                           n5143, ZN => n5893);
   U6321 : AOI22_X1 port map( A1 => n5786, A2 => n5144, B1 => n5787, B2 => 
                           n5145, ZN => n5892);
   U6322 : NAND3_X1 port map( A1 => n5896, A2 => n5897, A3 => n5898, ZN => 
                           n12996);
   U6323 : AOI221_X1 port map( B1 => n5779, B2 => n5149, C1 => n5780, C2 => 
                           MEM_IN(28), A => n5899, ZN => n5898);
   U6324 : OAI22_X1 port map( A1 => n11633, A2 => n235, B1 => n5151, B2 => 
                           n5783, ZN => n5899);
   U6325 : AOI22_X1 port map( A1 => n5784, A2 => n5152, B1 => n5785, B2 => 
                           n5153, ZN => n5897);
   U6326 : AOI22_X1 port map( A1 => n5786, A2 => n5154, B1 => n5787, B2 => 
                           n5155, ZN => n5896);
   U6327 : NAND3_X1 port map( A1 => n5900, A2 => n5901, A3 => n5902, ZN => 
                           n12995);
   U6328 : AOI221_X1 port map( B1 => n5779, B2 => n5159, C1 => n5780, C2 => 
                           MEM_IN(29), A => n5903, ZN => n5902);
   U6329 : OAI22_X1 port map( A1 => n11632, A2 => n235, B1 => n5161, B2 => 
                           n5783, ZN => n5903);
   U6330 : AOI22_X1 port map( A1 => n5784, A2 => n5162, B1 => n5785, B2 => 
                           n5163, ZN => n5901);
   U6331 : AOI22_X1 port map( A1 => n5786, A2 => n5164, B1 => n5787, B2 => 
                           n5165, ZN => n5900);
   U6332 : NAND3_X1 port map( A1 => n5904, A2 => n5905, A3 => n5906, ZN => 
                           n12994);
   U6333 : AOI221_X1 port map( B1 => n5779, B2 => n5169, C1 => n5780, C2 => 
                           MEM_IN(30), A => n5907, ZN => n5906);
   U6334 : OAI22_X1 port map( A1 => n11631, A2 => n235, B1 => n5171, B2 => 
                           n5783, ZN => n5907);
   U6335 : AOI22_X1 port map( A1 => n5784, A2 => n5172, B1 => n5785, B2 => 
                           n5173, ZN => n5905);
   U6336 : AOI22_X1 port map( A1 => n5786, A2 => n5174, B1 => n5787, B2 => 
                           n5175, ZN => n5904);
   U6337 : NAND3_X1 port map( A1 => n5908, A2 => n5909, A3 => n5910, ZN => 
                           n12993);
   U6338 : AOI221_X1 port map( B1 => n5779, B2 => n5179, C1 => n5780, C2 => 
                           MEM_IN(31), A => n5911, ZN => n5910);
   U6339 : OAI22_X1 port map( A1 => n11630, A2 => n235, B1 => n5181, B2 => 
                           n5783, ZN => n5911);
   U6340 : AOI22_X1 port map( A1 => n5784, A2 => n5191, B1 => n5785, B2 => 
                           n5192, ZN => n5909);
   U6341 : AOI22_X1 port map( A1 => n5786, A2 => n5195, B1 => n5787, B2 => 
                           n5196, ZN => n5908);
   U6342 : OAI22_X1 port map( A1 => n5914, A2 => n5919, B1 => n208, B2 => n234,
                           ZN => n5915);
   U6343 : INV_X1 port map( A => n5913, ZN => n5919);
   U6344 : NOR3_X1 port map( A1 => n4841, A2 => n234, A3 => n5912, ZN => n5913)
                           ;
   U6345 : OAI22_X1 port map( A1 => n4786, A2 => n5920, B1 => n5921, B2 => 
                           n5204, ZN => n5782);
   U6346 : NOR2_X1 port map( A1 => n5914, A2 => n5912, ZN => n5921);
   U6347 : NAND4_X1 port map( A1 => n5767, A2 => n5516, A3 => n5772, A4 => 
                           n5774, ZN => n5912);
   U6348 : NOR4_X1 port map( A1 => n5922, A2 => n5769, A3 => RESET, A4 => n5917
                           , ZN => n5920);
   U6349 : OAI211_X1 port map( C1 => n5770, C2 => n5923, A => n5756, B => n5515
                           , ZN => n5922);
   U6350 : INV_X1 port map( A => n5517, ZN => n5515);
   U6351 : INV_X1 port map( A => n5360, ZN => n5756);
   U6352 : NOR2_X1 port map( A1 => n5516, A2 => n4787, ZN => n5360);
   U6353 : NAND2_X1 port map( A1 => n5924, A2 => n5925, ZN => n5914);
   U6354 : INV_X1 port map( A => n5516, ZN => n5359);
   U6355 : NAND2_X1 port map( A1 => n5926, A2 => n5216, ZN => n5516);
   U6356 : NAND3_X1 port map( A1 => n5927, A2 => n5928, A3 => n5929, ZN => 
                           n12992);
   U6357 : AOI221_X1 port map( B1 => n5930, B2 => n4863, C1 => n5931, C2 => 
                           MEM_IN(0), A => n5932, ZN => n5929);
   U6358 : OAI22_X1 port map( A1 => n11629, A2 => n222, B1 => n4867, B2 => 
                           n5934, ZN => n5932);
   U6359 : AOI22_X1 port map( A1 => n5935, A2 => n4869, B1 => n5936, B2 => 
                           n4871, ZN => n5928);
   U6360 : AOI22_X1 port map( A1 => n5937, A2 => n4873, B1 => n5938, B2 => 
                           n4875, ZN => n5927);
   U6361 : NAND3_X1 port map( A1 => n5939, A2 => n5940, A3 => n5941, ZN => 
                           n12991);
   U6362 : AOI221_X1 port map( B1 => n5930, B2 => n4879, C1 => n5931, C2 => 
                           MEM_IN(1), A => n5942, ZN => n5941);
   U6363 : OAI22_X1 port map( A1 => n11628, A2 => n222, B1 => n4881, B2 => 
                           n5934, ZN => n5942);
   U6364 : AOI22_X1 port map( A1 => n5935, A2 => n4882, B1 => n5936, B2 => 
                           n4883, ZN => n5940);
   U6365 : AOI22_X1 port map( A1 => n5937, A2 => n4884, B1 => n5938, B2 => 
                           n4885, ZN => n5939);
   U6366 : NAND3_X1 port map( A1 => n5943, A2 => n5944, A3 => n5945, ZN => 
                           n12990);
   U6367 : AOI221_X1 port map( B1 => n5930, B2 => n4889, C1 => n5931, C2 => 
                           MEM_IN(2), A => n5946, ZN => n5945);
   U6368 : OAI22_X1 port map( A1 => n11627, A2 => n222, B1 => n4891, B2 => 
                           n5934, ZN => n5946);
   U6369 : AOI22_X1 port map( A1 => n5935, A2 => n4892, B1 => n5936, B2 => 
                           n4893, ZN => n5944);
   U6370 : AOI22_X1 port map( A1 => n5937, A2 => n4894, B1 => n5938, B2 => 
                           n4895, ZN => n5943);
   U6371 : NAND3_X1 port map( A1 => n5947, A2 => n5948, A3 => n5949, ZN => 
                           n12989);
   U6372 : AOI221_X1 port map( B1 => n5930, B2 => n4899, C1 => n5931, C2 => 
                           MEM_IN(3), A => n5950, ZN => n5949);
   U6373 : OAI22_X1 port map( A1 => n11626, A2 => n222, B1 => n4901, B2 => 
                           n5934, ZN => n5950);
   U6374 : AOI22_X1 port map( A1 => n5935, A2 => n4902, B1 => n5936, B2 => 
                           n4903, ZN => n5948);
   U6375 : AOI22_X1 port map( A1 => n5937, A2 => n4904, B1 => n5938, B2 => 
                           n4905, ZN => n5947);
   U6376 : NAND3_X1 port map( A1 => n5951, A2 => n5952, A3 => n5953, ZN => 
                           n12988);
   U6377 : AOI221_X1 port map( B1 => n5930, B2 => n4909, C1 => n5931, C2 => 
                           MEM_IN(4), A => n5954, ZN => n5953);
   U6378 : OAI22_X1 port map( A1 => n11625, A2 => n222, B1 => n4911, B2 => 
                           n5934, ZN => n5954);
   U6379 : AOI22_X1 port map( A1 => n5935, A2 => n4912, B1 => n5936, B2 => 
                           n4913, ZN => n5952);
   U6380 : AOI22_X1 port map( A1 => n5937, A2 => n4914, B1 => n5938, B2 => 
                           n4915, ZN => n5951);
   U6381 : NAND3_X1 port map( A1 => n5955, A2 => n5956, A3 => n5957, ZN => 
                           n12987);
   U6382 : AOI221_X1 port map( B1 => n5930, B2 => n4919, C1 => n5931, C2 => 
                           MEM_IN(5), A => n5958, ZN => n5957);
   U6383 : OAI22_X1 port map( A1 => n11624, A2 => n222, B1 => n4921, B2 => 
                           n5934, ZN => n5958);
   U6384 : AOI22_X1 port map( A1 => n5935, A2 => n4922, B1 => n5936, B2 => 
                           n4923, ZN => n5956);
   U6385 : AOI22_X1 port map( A1 => n5937, A2 => n4924, B1 => n5938, B2 => 
                           n4925, ZN => n5955);
   U6386 : NAND3_X1 port map( A1 => n5959, A2 => n5960, A3 => n5961, ZN => 
                           n12986);
   U6387 : AOI221_X1 port map( B1 => n5930, B2 => n4929, C1 => n5931, C2 => 
                           MEM_IN(6), A => n5962, ZN => n5961);
   U6388 : OAI22_X1 port map( A1 => n11623, A2 => n222, B1 => n4931, B2 => 
                           n5934, ZN => n5962);
   U6389 : AOI22_X1 port map( A1 => n5935, A2 => n4932, B1 => n5936, B2 => 
                           n4933, ZN => n5960);
   U6390 : AOI22_X1 port map( A1 => n5937, A2 => n4934, B1 => n5938, B2 => 
                           n4935, ZN => n5959);
   U6391 : NAND3_X1 port map( A1 => n5963, A2 => n5964, A3 => n5965, ZN => 
                           n12985);
   U6392 : AOI221_X1 port map( B1 => n5930, B2 => n4939, C1 => n5931, C2 => 
                           MEM_IN(7), A => n5966, ZN => n5965);
   U6393 : OAI22_X1 port map( A1 => n11622, A2 => n222, B1 => n4941, B2 => 
                           n5934, ZN => n5966);
   U6394 : AOI22_X1 port map( A1 => n5935, A2 => n4942, B1 => n5936, B2 => 
                           n4943, ZN => n5964);
   U6395 : AOI22_X1 port map( A1 => n5937, A2 => n4944, B1 => n5938, B2 => 
                           n4945, ZN => n5963);
   U6396 : NAND3_X1 port map( A1 => n5967, A2 => n5968, A3 => n5969, ZN => 
                           n12984);
   U6397 : AOI221_X1 port map( B1 => n5930, B2 => n4949, C1 => n5931, C2 => 
                           MEM_IN(8), A => n5970, ZN => n5969);
   U6398 : OAI22_X1 port map( A1 => n11621, A2 => n222, B1 => n4951, B2 => 
                           n5934, ZN => n5970);
   U6399 : AOI22_X1 port map( A1 => n5935, A2 => n4952, B1 => n5936, B2 => 
                           n4953, ZN => n5968);
   U6400 : AOI22_X1 port map( A1 => n5937, A2 => n4954, B1 => n5938, B2 => 
                           n4955, ZN => n5967);
   U6401 : NAND3_X1 port map( A1 => n5971, A2 => n5972, A3 => n5973, ZN => 
                           n12983);
   U6402 : AOI221_X1 port map( B1 => n5930, B2 => n4959, C1 => n5931, C2 => 
                           MEM_IN(9), A => n5974, ZN => n5973);
   U6403 : OAI22_X1 port map( A1 => n11620, A2 => n222, B1 => n4961, B2 => 
                           n5934, ZN => n5974);
   U6404 : AOI22_X1 port map( A1 => n5935, A2 => n4962, B1 => n5936, B2 => 
                           n4963, ZN => n5972);
   U6405 : AOI22_X1 port map( A1 => n5937, A2 => n4964, B1 => n5938, B2 => 
                           n4965, ZN => n5971);
   U6406 : NAND3_X1 port map( A1 => n5975, A2 => n5976, A3 => n5977, ZN => 
                           n12982);
   U6407 : AOI221_X1 port map( B1 => n5930, B2 => n4969, C1 => n5931, C2 => 
                           MEM_IN(10), A => n5978, ZN => n5977);
   U6408 : OAI22_X1 port map( A1 => n11619, A2 => n222, B1 => n4971, B2 => 
                           n5934, ZN => n5978);
   U6409 : AOI22_X1 port map( A1 => n5935, A2 => n4972, B1 => n5936, B2 => 
                           n4973, ZN => n5976);
   U6410 : AOI22_X1 port map( A1 => n5937, A2 => n4974, B1 => n5938, B2 => 
                           n4975, ZN => n5975);
   U6411 : NAND3_X1 port map( A1 => n5979, A2 => n5980, A3 => n5981, ZN => 
                           n12981);
   U6412 : AOI221_X1 port map( B1 => n5930, B2 => n4979, C1 => n5931, C2 => 
                           MEM_IN(11), A => n5982, ZN => n5981);
   U6413 : OAI22_X1 port map( A1 => n11618, A2 => n222, B1 => n4981, B2 => 
                           n5934, ZN => n5982);
   U6414 : AOI22_X1 port map( A1 => n5935, A2 => n4982, B1 => n5936, B2 => 
                           n4983, ZN => n5980);
   U6415 : AOI22_X1 port map( A1 => n5937, A2 => n4984, B1 => n5938, B2 => 
                           n4985, ZN => n5979);
   U6416 : NAND3_X1 port map( A1 => n5983, A2 => n5984, A3 => n5985, ZN => 
                           n12980);
   U6417 : AOI221_X1 port map( B1 => n5930, B2 => n4989, C1 => n5931, C2 => 
                           MEM_IN(12), A => n5986, ZN => n5985);
   U6418 : OAI22_X1 port map( A1 => n11617, A2 => n222, B1 => n4991, B2 => 
                           n5934, ZN => n5986);
   U6419 : AOI22_X1 port map( A1 => n5935, A2 => n4992, B1 => n5936, B2 => 
                           n4993, ZN => n5984);
   U6420 : AOI22_X1 port map( A1 => n5937, A2 => n4994, B1 => n5938, B2 => 
                           n4995, ZN => n5983);
   U6421 : NAND3_X1 port map( A1 => n5987, A2 => n5988, A3 => n5989, ZN => 
                           n12979);
   U6422 : AOI221_X1 port map( B1 => n5930, B2 => n4999, C1 => n5931, C2 => 
                           MEM_IN(13), A => n5990, ZN => n5989);
   U6423 : OAI22_X1 port map( A1 => n11616, A2 => n222, B1 => n5001, B2 => 
                           n5934, ZN => n5990);
   U6424 : AOI22_X1 port map( A1 => n5935, A2 => n5002, B1 => n5936, B2 => 
                           n5003, ZN => n5988);
   U6425 : AOI22_X1 port map( A1 => n5937, A2 => n5004, B1 => n5938, B2 => 
                           n5005, ZN => n5987);
   U6426 : NAND3_X1 port map( A1 => n5991, A2 => n5992, A3 => n5993, ZN => 
                           n12978);
   U6427 : AOI221_X1 port map( B1 => n5930, B2 => n5009, C1 => n5931, C2 => 
                           MEM_IN(14), A => n5994, ZN => n5993);
   U6428 : OAI22_X1 port map( A1 => n11615, A2 => n222, B1 => n5011, B2 => 
                           n5934, ZN => n5994);
   U6429 : AOI22_X1 port map( A1 => n5935, A2 => n5012, B1 => n5936, B2 => 
                           n5013, ZN => n5992);
   U6430 : AOI22_X1 port map( A1 => n5937, A2 => n5014, B1 => n5938, B2 => 
                           n5015, ZN => n5991);
   U6431 : NAND3_X1 port map( A1 => n5995, A2 => n5996, A3 => n5997, ZN => 
                           n12977);
   U6432 : AOI221_X1 port map( B1 => n5930, B2 => n5019, C1 => n5931, C2 => 
                           MEM_IN(15), A => n5998, ZN => n5997);
   U6433 : OAI22_X1 port map( A1 => n11614, A2 => n222, B1 => n5021, B2 => 
                           n5934, ZN => n5998);
   U6434 : AOI22_X1 port map( A1 => n5935, A2 => n5022, B1 => n5936, B2 => 
                           n5023, ZN => n5996);
   U6435 : AOI22_X1 port map( A1 => n5937, A2 => n5024, B1 => n5938, B2 => 
                           n5025, ZN => n5995);
   U6436 : NAND3_X1 port map( A1 => n5999, A2 => n6000, A3 => n6001, ZN => 
                           n12976);
   U6437 : AOI221_X1 port map( B1 => n5930, B2 => n5029, C1 => n5931, C2 => 
                           MEM_IN(16), A => n6002, ZN => n6001);
   U6438 : OAI22_X1 port map( A1 => n11613, A2 => n222, B1 => n5031, B2 => 
                           n5934, ZN => n6002);
   U6439 : AOI22_X1 port map( A1 => n5935, A2 => n5032, B1 => n5936, B2 => 
                           n5033, ZN => n6000);
   U6440 : AOI22_X1 port map( A1 => n5937, A2 => n5034, B1 => n5938, B2 => 
                           n5035, ZN => n5999);
   U6441 : NAND3_X1 port map( A1 => n6003, A2 => n6004, A3 => n6005, ZN => 
                           n12975);
   U6442 : AOI221_X1 port map( B1 => n5930, B2 => n5039, C1 => n5931, C2 => 
                           MEM_IN(17), A => n6006, ZN => n6005);
   U6443 : OAI22_X1 port map( A1 => n11612, A2 => n222, B1 => n5041, B2 => 
                           n5934, ZN => n6006);
   U6444 : AOI22_X1 port map( A1 => n5935, A2 => n5042, B1 => n5936, B2 => 
                           n5043, ZN => n6004);
   U6445 : AOI22_X1 port map( A1 => n5937, A2 => n5044, B1 => n5938, B2 => 
                           n5045, ZN => n6003);
   U6446 : NAND3_X1 port map( A1 => n6007, A2 => n6008, A3 => n6009, ZN => 
                           n12974);
   U6447 : AOI221_X1 port map( B1 => n5930, B2 => n5049, C1 => n5931, C2 => 
                           MEM_IN(18), A => n6010, ZN => n6009);
   U6448 : OAI22_X1 port map( A1 => n11611, A2 => n222, B1 => n5051, B2 => 
                           n5934, ZN => n6010);
   U6449 : AOI22_X1 port map( A1 => n5935, A2 => n5052, B1 => n5936, B2 => 
                           n5053, ZN => n6008);
   U6450 : AOI22_X1 port map( A1 => n5937, A2 => n5054, B1 => n5938, B2 => 
                           n5055, ZN => n6007);
   U6451 : NAND3_X1 port map( A1 => n6011, A2 => n6012, A3 => n6013, ZN => 
                           n12973);
   U6452 : AOI221_X1 port map( B1 => n5930, B2 => n5059, C1 => n5931, C2 => 
                           MEM_IN(19), A => n6014, ZN => n6013);
   U6453 : OAI22_X1 port map( A1 => n11610, A2 => n222, B1 => n5061, B2 => 
                           n5934, ZN => n6014);
   U6454 : AOI22_X1 port map( A1 => n5935, A2 => n5062, B1 => n5936, B2 => 
                           n5063, ZN => n6012);
   U6455 : AOI22_X1 port map( A1 => n5937, A2 => n5064, B1 => n5938, B2 => 
                           n5065, ZN => n6011);
   U6456 : NAND3_X1 port map( A1 => n6015, A2 => n6016, A3 => n6017, ZN => 
                           n12972);
   U6457 : AOI221_X1 port map( B1 => n5930, B2 => n5069, C1 => n5931, C2 => 
                           MEM_IN(20), A => n6018, ZN => n6017);
   U6458 : OAI22_X1 port map( A1 => n11609, A2 => n222, B1 => n5071, B2 => 
                           n5934, ZN => n6018);
   U6459 : AOI22_X1 port map( A1 => n5935, A2 => n5072, B1 => n5936, B2 => 
                           n5073, ZN => n6016);
   U6460 : AOI22_X1 port map( A1 => n5937, A2 => n5074, B1 => n5938, B2 => 
                           n5075, ZN => n6015);
   U6461 : NAND3_X1 port map( A1 => n6019, A2 => n6020, A3 => n6021, ZN => 
                           n12971);
   U6462 : AOI221_X1 port map( B1 => n5930, B2 => n5079, C1 => n5931, C2 => 
                           MEM_IN(21), A => n6022, ZN => n6021);
   U6463 : OAI22_X1 port map( A1 => n11608, A2 => n222, B1 => n5081, B2 => 
                           n5934, ZN => n6022);
   U6464 : AOI22_X1 port map( A1 => n5935, A2 => n5082, B1 => n5936, B2 => 
                           n5083, ZN => n6020);
   U6465 : AOI22_X1 port map( A1 => n5937, A2 => n5084, B1 => n5938, B2 => 
                           n5085, ZN => n6019);
   U6466 : NAND3_X1 port map( A1 => n6023, A2 => n6024, A3 => n6025, ZN => 
                           n12970);
   U6467 : AOI221_X1 port map( B1 => n5930, B2 => n5089, C1 => n5931, C2 => 
                           MEM_IN(22), A => n6026, ZN => n6025);
   U6468 : OAI22_X1 port map( A1 => n11607, A2 => n222, B1 => n5091, B2 => 
                           n5934, ZN => n6026);
   U6469 : AOI22_X1 port map( A1 => n5935, A2 => n5092, B1 => n5936, B2 => 
                           n5093, ZN => n6024);
   U6470 : AOI22_X1 port map( A1 => n5937, A2 => n5094, B1 => n5938, B2 => 
                           n5095, ZN => n6023);
   U6471 : NAND3_X1 port map( A1 => n6027, A2 => n6028, A3 => n6029, ZN => 
                           n12969);
   U6472 : AOI221_X1 port map( B1 => n5930, B2 => n5099, C1 => n5931, C2 => 
                           MEM_IN(23), A => n6030, ZN => n6029);
   U6473 : OAI22_X1 port map( A1 => n11606, A2 => n222, B1 => n5101, B2 => 
                           n5934, ZN => n6030);
   U6474 : AOI22_X1 port map( A1 => n5935, A2 => n5102, B1 => n5936, B2 => 
                           n5103, ZN => n6028);
   U6475 : AOI22_X1 port map( A1 => n5937, A2 => n5104, B1 => n5938, B2 => 
                           n5105, ZN => n6027);
   U6476 : NAND3_X1 port map( A1 => n6031, A2 => n6032, A3 => n6033, ZN => 
                           n12968);
   U6477 : AOI221_X1 port map( B1 => n5930, B2 => n5109, C1 => n5931, C2 => 
                           MEM_IN(24), A => n6034, ZN => n6033);
   U6478 : OAI22_X1 port map( A1 => n11605, A2 => n222, B1 => n5111, B2 => 
                           n5934, ZN => n6034);
   U6479 : AOI22_X1 port map( A1 => n5935, A2 => n5112, B1 => n5936, B2 => 
                           n5113, ZN => n6032);
   U6480 : AOI22_X1 port map( A1 => n5937, A2 => n5114, B1 => n5938, B2 => 
                           n5115, ZN => n6031);
   U6481 : NAND3_X1 port map( A1 => n6035, A2 => n6036, A3 => n6037, ZN => 
                           n12967);
   U6482 : AOI221_X1 port map( B1 => n5930, B2 => n5119, C1 => n5931, C2 => 
                           MEM_IN(25), A => n6038, ZN => n6037);
   U6483 : OAI22_X1 port map( A1 => n11604, A2 => n222, B1 => n5121, B2 => 
                           n5934, ZN => n6038);
   U6484 : AOI22_X1 port map( A1 => n5935, A2 => n5122, B1 => n5936, B2 => 
                           n5123, ZN => n6036);
   U6485 : AOI22_X1 port map( A1 => n5937, A2 => n5124, B1 => n5938, B2 => 
                           n5125, ZN => n6035);
   U6486 : NAND3_X1 port map( A1 => n6039, A2 => n6040, A3 => n6041, ZN => 
                           n12966);
   U6487 : AOI221_X1 port map( B1 => n5930, B2 => n5129, C1 => n5931, C2 => 
                           MEM_IN(26), A => n6042, ZN => n6041);
   U6488 : OAI22_X1 port map( A1 => n11603, A2 => n222, B1 => n5131, B2 => 
                           n5934, ZN => n6042);
   U6489 : AOI22_X1 port map( A1 => n5935, A2 => n5132, B1 => n5936, B2 => 
                           n5133, ZN => n6040);
   U6490 : AOI22_X1 port map( A1 => n5937, A2 => n5134, B1 => n5938, B2 => 
                           n5135, ZN => n6039);
   U6491 : NAND3_X1 port map( A1 => n6043, A2 => n6044, A3 => n6045, ZN => 
                           n12965);
   U6492 : AOI221_X1 port map( B1 => n5930, B2 => n5139, C1 => n5931, C2 => 
                           MEM_IN(27), A => n6046, ZN => n6045);
   U6493 : OAI22_X1 port map( A1 => n11602, A2 => n222, B1 => n5141, B2 => 
                           n5934, ZN => n6046);
   U6494 : AOI22_X1 port map( A1 => n5935, A2 => n5142, B1 => n5936, B2 => 
                           n5143, ZN => n6044);
   U6495 : AOI22_X1 port map( A1 => n5937, A2 => n5144, B1 => n5938, B2 => 
                           n5145, ZN => n6043);
   U6496 : NAND3_X1 port map( A1 => n6047, A2 => n6048, A3 => n6049, ZN => 
                           n12964);
   U6497 : AOI221_X1 port map( B1 => n5930, B2 => n5149, C1 => n5931, C2 => 
                           MEM_IN(28), A => n6050, ZN => n6049);
   U6498 : OAI22_X1 port map( A1 => n11601, A2 => n222, B1 => n5151, B2 => 
                           n5934, ZN => n6050);
   U6499 : AOI22_X1 port map( A1 => n5935, A2 => n5152, B1 => n5936, B2 => 
                           n5153, ZN => n6048);
   U6500 : AOI22_X1 port map( A1 => n5937, A2 => n5154, B1 => n5938, B2 => 
                           n5155, ZN => n6047);
   U6501 : NAND3_X1 port map( A1 => n6051, A2 => n6052, A3 => n6053, ZN => 
                           n12963);
   U6502 : AOI221_X1 port map( B1 => n5930, B2 => n5159, C1 => n5931, C2 => 
                           MEM_IN(29), A => n6054, ZN => n6053);
   U6503 : OAI22_X1 port map( A1 => n11600, A2 => n222, B1 => n5161, B2 => 
                           n5934, ZN => n6054);
   U6504 : AOI22_X1 port map( A1 => n5935, A2 => n5162, B1 => n5936, B2 => 
                           n5163, ZN => n6052);
   U6505 : AOI22_X1 port map( A1 => n5937, A2 => n5164, B1 => n5938, B2 => 
                           n5165, ZN => n6051);
   U6506 : NAND3_X1 port map( A1 => n6055, A2 => n6056, A3 => n6057, ZN => 
                           n12962);
   U6507 : AOI221_X1 port map( B1 => n5930, B2 => n5169, C1 => n5931, C2 => 
                           MEM_IN(30), A => n6058, ZN => n6057);
   U6508 : OAI22_X1 port map( A1 => n11599, A2 => n222, B1 => n5171, B2 => 
                           n5934, ZN => n6058);
   U6509 : AOI22_X1 port map( A1 => n5935, A2 => n5172, B1 => n5936, B2 => 
                           n5173, ZN => n6056);
   U6510 : AOI22_X1 port map( A1 => n5937, A2 => n5174, B1 => n5938, B2 => 
                           n5175, ZN => n6055);
   U6511 : NAND3_X1 port map( A1 => n6059, A2 => n6060, A3 => n6061, ZN => 
                           n12961);
   U6512 : AOI221_X1 port map( B1 => n5930, B2 => n5179, C1 => n5931, C2 => 
                           MEM_IN(31), A => n6062, ZN => n6061);
   U6513 : OAI22_X1 port map( A1 => n11598, A2 => n222, B1 => n5181, B2 => 
                           n5934, ZN => n6062);
   U6514 : OR2_X1 port map( A1 => n4787, A2 => n5918, ZN => n5916);
   U6515 : AND4_X1 port map( A1 => n5206, A2 => n5772, A3 => n6068, A4 => n5521
                           , ZN => n5918);
   U6516 : AOI22_X1 port map( A1 => n5935, A2 => n5191, B1 => n5936, B2 => 
                           n5192, ZN => n6060);
   U6517 : AOI22_X1 port map( A1 => n5937, A2 => n5195, B1 => n5938, B2 => 
                           n5196, ZN => n6059);
   U6518 : OAI22_X1 port map( A1 => n6065, A2 => n6070, B1 => n208, B2 => n221,
                           ZN => n6067);
   U6519 : INV_X1 port map( A => n6064, ZN => n6070);
   U6520 : NOR3_X1 port map( A1 => n4841, A2 => n221, A3 => n6063, ZN => n6064)
                           ;
   U6521 : OAI22_X1 port map( A1 => n4786, A2 => n6071, B1 => n6072, B2 => 
                           n5204, ZN => n5933);
   U6522 : NOR2_X1 port map( A1 => n6065, A2 => n6063, ZN => n6072);
   U6523 : NAND3_X1 port map( A1 => n6073, A2 => n5772, A3 => n5767, ZN => 
                           n6063);
   U6524 : INV_X1 port map( A => n6074, ZN => n6073);
   U6525 : NOR3_X1 port map( A1 => n6075, A2 => RESET, A3 => n5517, ZN => n6071
                           );
   U6526 : OAI22_X1 port map( A1 => n5770, A2 => n6076, B1 => n5767, B2 => 
                           n4787, ZN => n6075);
   U6527 : OR2_X1 port map( A1 => n6077, A2 => n6078, ZN => n6065);
   U6528 : NOR2_X1 port map( A1 => n5772, A2 => n4787, ZN => n5517);
   U6529 : NAND2_X1 port map( A1 => n6079, A2 => n5216, ZN => n5772);
   U6530 : NAND3_X1 port map( A1 => n6080, A2 => n6081, A3 => n6082, ZN => 
                           n12960);
   U6531 : AOI221_X1 port map( B1 => n151, B2 => n4863, C1 => n6083, C2 => 
                           MEM_IN(0), A => n6084, ZN => n6082);
   U6532 : OAI22_X1 port map( A1 => n11597, A2 => n6085, B1 => n4867, B2 => 
                           n6086, ZN => n6084);
   U6533 : AOI22_X1 port map( A1 => n204, A2 => n4869, B1 => n165, B2 => n4871,
                           ZN => n6081);
   U6534 : AOI22_X1 port map( A1 => n205, A2 => n4873, B1 => n162, B2 => n4875,
                           ZN => n6080);
   U6535 : NAND3_X1 port map( A1 => n6087, A2 => n6088, A3 => n6089, ZN => 
                           n12959);
   U6536 : AOI221_X1 port map( B1 => n151, B2 => n4879, C1 => n6083, C2 => 
                           MEM_IN(1), A => n6090, ZN => n6089);
   U6537 : OAI22_X1 port map( A1 => n11596, A2 => n6085, B1 => n4881, B2 => 
                           n6086, ZN => n6090);
   U6538 : AOI22_X1 port map( A1 => n204, A2 => n4882, B1 => n165, B2 => n4883,
                           ZN => n6088);
   U6539 : AOI22_X1 port map( A1 => n205, A2 => n4884, B1 => n162, B2 => n4885,
                           ZN => n6087);
   U6540 : NAND3_X1 port map( A1 => n6091, A2 => n6092, A3 => n6093, ZN => 
                           n12958);
   U6541 : AOI221_X1 port map( B1 => n151, B2 => n4889, C1 => n6083, C2 => 
                           MEM_IN(2), A => n6094, ZN => n6093);
   U6542 : OAI22_X1 port map( A1 => n11595, A2 => n6085, B1 => n4891, B2 => 
                           n6086, ZN => n6094);
   U6543 : AOI22_X1 port map( A1 => n204, A2 => n4892, B1 => n165, B2 => n4893,
                           ZN => n6092);
   U6544 : AOI22_X1 port map( A1 => n205, A2 => n4894, B1 => n162, B2 => n4895,
                           ZN => n6091);
   U6545 : NAND3_X1 port map( A1 => n6095, A2 => n6096, A3 => n6097, ZN => 
                           n12957);
   U6546 : AOI221_X1 port map( B1 => n151, B2 => n4899, C1 => n6083, C2 => 
                           MEM_IN(3), A => n6098, ZN => n6097);
   U6547 : OAI22_X1 port map( A1 => n11594, A2 => n6085, B1 => n4901, B2 => 
                           n6086, ZN => n6098);
   U6548 : AOI22_X1 port map( A1 => n204, A2 => n4902, B1 => n165, B2 => n4903,
                           ZN => n6096);
   U6549 : AOI22_X1 port map( A1 => n205, A2 => n4904, B1 => n162, B2 => n4905,
                           ZN => n6095);
   U6550 : NAND3_X1 port map( A1 => n6099, A2 => n6100, A3 => n6101, ZN => 
                           n12956);
   U6551 : AOI221_X1 port map( B1 => n151, B2 => n4909, C1 => n6083, C2 => 
                           MEM_IN(4), A => n6102, ZN => n6101);
   U6552 : OAI22_X1 port map( A1 => n11593, A2 => n6085, B1 => n4911, B2 => 
                           n6086, ZN => n6102);
   U6553 : AOI22_X1 port map( A1 => n204, A2 => n4912, B1 => n165, B2 => n4913,
                           ZN => n6100);
   U6554 : AOI22_X1 port map( A1 => n205, A2 => n4914, B1 => n162, B2 => n4915,
                           ZN => n6099);
   U6555 : NAND3_X1 port map( A1 => n6103, A2 => n6104, A3 => n6105, ZN => 
                           n12955);
   U6556 : AOI221_X1 port map( B1 => n151, B2 => n4919, C1 => n6083, C2 => 
                           MEM_IN(5), A => n6106, ZN => n6105);
   U6557 : OAI22_X1 port map( A1 => n11592, A2 => n6085, B1 => n4921, B2 => 
                           n6086, ZN => n6106);
   U6558 : AOI22_X1 port map( A1 => n204, A2 => n4922, B1 => n165, B2 => n4923,
                           ZN => n6104);
   U6559 : AOI22_X1 port map( A1 => n205, A2 => n4924, B1 => n162, B2 => n4925,
                           ZN => n6103);
   U6560 : NAND3_X1 port map( A1 => n6107, A2 => n6108, A3 => n6109, ZN => 
                           n12954);
   U6561 : AOI221_X1 port map( B1 => n151, B2 => n4929, C1 => n6083, C2 => 
                           MEM_IN(6), A => n6110, ZN => n6109);
   U6562 : OAI22_X1 port map( A1 => n11591, A2 => n6085, B1 => n4931, B2 => 
                           n6086, ZN => n6110);
   U6563 : AOI22_X1 port map( A1 => n204, A2 => n4932, B1 => n165, B2 => n4933,
                           ZN => n6108);
   U6564 : AOI22_X1 port map( A1 => n205, A2 => n4934, B1 => n162, B2 => n4935,
                           ZN => n6107);
   U6565 : NAND3_X1 port map( A1 => n6111, A2 => n6112, A3 => n6113, ZN => 
                           n12953);
   U6566 : AOI221_X1 port map( B1 => n151, B2 => n4939, C1 => n6083, C2 => 
                           MEM_IN(7), A => n6114, ZN => n6113);
   U6567 : OAI22_X1 port map( A1 => n11590, A2 => n6085, B1 => n4941, B2 => 
                           n6086, ZN => n6114);
   U6568 : AOI22_X1 port map( A1 => n204, A2 => n4942, B1 => n165, B2 => n4943,
                           ZN => n6112);
   U6569 : AOI22_X1 port map( A1 => n205, A2 => n4944, B1 => n162, B2 => n4945,
                           ZN => n6111);
   U6570 : NAND3_X1 port map( A1 => n6115, A2 => n6116, A3 => n6117, ZN => 
                           n12952);
   U6571 : AOI221_X1 port map( B1 => n151, B2 => n4949, C1 => n6083, C2 => 
                           MEM_IN(8), A => n6118, ZN => n6117);
   U6572 : OAI22_X1 port map( A1 => n11589, A2 => n6085, B1 => n4951, B2 => 
                           n6086, ZN => n6118);
   U6573 : AOI22_X1 port map( A1 => n204, A2 => n4952, B1 => n165, B2 => n4953,
                           ZN => n6116);
   U6574 : AOI22_X1 port map( A1 => n205, A2 => n4954, B1 => n162, B2 => n4955,
                           ZN => n6115);
   U6575 : NAND3_X1 port map( A1 => n6119, A2 => n6120, A3 => n6121, ZN => 
                           n12951);
   U6576 : AOI221_X1 port map( B1 => n151, B2 => n4959, C1 => n6083, C2 => 
                           MEM_IN(9), A => n6122, ZN => n6121);
   U6577 : OAI22_X1 port map( A1 => n11588, A2 => n6085, B1 => n4961, B2 => 
                           n6086, ZN => n6122);
   U6578 : AOI22_X1 port map( A1 => n204, A2 => n4962, B1 => n165, B2 => n4963,
                           ZN => n6120);
   U6579 : AOI22_X1 port map( A1 => n205, A2 => n4964, B1 => n162, B2 => n4965,
                           ZN => n6119);
   U6580 : NAND3_X1 port map( A1 => n6123, A2 => n6124, A3 => n6125, ZN => 
                           n12950);
   U6581 : AOI221_X1 port map( B1 => n151, B2 => n4969, C1 => n6083, C2 => 
                           MEM_IN(10), A => n6126, ZN => n6125);
   U6582 : OAI22_X1 port map( A1 => n11587, A2 => n6085, B1 => n4971, B2 => 
                           n6086, ZN => n6126);
   U6583 : AOI22_X1 port map( A1 => n204, A2 => n4972, B1 => n165, B2 => n4973,
                           ZN => n6124);
   U6584 : AOI22_X1 port map( A1 => n205, A2 => n4974, B1 => n162, B2 => n4975,
                           ZN => n6123);
   U6585 : NAND3_X1 port map( A1 => n6127, A2 => n6128, A3 => n6129, ZN => 
                           n12949);
   U6586 : AOI221_X1 port map( B1 => n151, B2 => n4979, C1 => n6083, C2 => 
                           MEM_IN(11), A => n6130, ZN => n6129);
   U6587 : OAI22_X1 port map( A1 => n11586, A2 => n6085, B1 => n4981, B2 => 
                           n6086, ZN => n6130);
   U6588 : AOI22_X1 port map( A1 => n204, A2 => n4982, B1 => n165, B2 => n4983,
                           ZN => n6128);
   U6589 : AOI22_X1 port map( A1 => n205, A2 => n4984, B1 => n162, B2 => n4985,
                           ZN => n6127);
   U6590 : NAND3_X1 port map( A1 => n6131, A2 => n6132, A3 => n6133, ZN => 
                           n12948);
   U6591 : AOI221_X1 port map( B1 => n151, B2 => n4989, C1 => n6083, C2 => 
                           MEM_IN(12), A => n6134, ZN => n6133);
   U6592 : OAI22_X1 port map( A1 => n11585, A2 => n6085, B1 => n4991, B2 => 
                           n6086, ZN => n6134);
   U6593 : AOI22_X1 port map( A1 => n204, A2 => n4992, B1 => n165, B2 => n4993,
                           ZN => n6132);
   U6594 : AOI22_X1 port map( A1 => n205, A2 => n4994, B1 => n162, B2 => n4995,
                           ZN => n6131);
   U6595 : NAND3_X1 port map( A1 => n6135, A2 => n6136, A3 => n6137, ZN => 
                           n12947);
   U6596 : AOI221_X1 port map( B1 => n151, B2 => n4999, C1 => n6083, C2 => 
                           MEM_IN(13), A => n6138, ZN => n6137);
   U6597 : OAI22_X1 port map( A1 => n11584, A2 => n6085, B1 => n5001, B2 => 
                           n6086, ZN => n6138);
   U6598 : AOI22_X1 port map( A1 => n204, A2 => n5002, B1 => n165, B2 => n5003,
                           ZN => n6136);
   U6599 : AOI22_X1 port map( A1 => n205, A2 => n5004, B1 => n162, B2 => n5005,
                           ZN => n6135);
   U6600 : NAND3_X1 port map( A1 => n6139, A2 => n6140, A3 => n6141, ZN => 
                           n12946);
   U6601 : AOI221_X1 port map( B1 => n151, B2 => n5009, C1 => n6083, C2 => 
                           MEM_IN(14), A => n6142, ZN => n6141);
   U6602 : OAI22_X1 port map( A1 => n11583, A2 => n6085, B1 => n5011, B2 => 
                           n6086, ZN => n6142);
   U6603 : AOI22_X1 port map( A1 => n204, A2 => n5012, B1 => n165, B2 => n5013,
                           ZN => n6140);
   U6604 : AOI22_X1 port map( A1 => n205, A2 => n5014, B1 => n162, B2 => n5015,
                           ZN => n6139);
   U6605 : NAND3_X1 port map( A1 => n6143, A2 => n6144, A3 => n6145, ZN => 
                           n12945);
   U6606 : AOI221_X1 port map( B1 => n151, B2 => n5019, C1 => n6083, C2 => 
                           MEM_IN(15), A => n6146, ZN => n6145);
   U6607 : OAI22_X1 port map( A1 => n11582, A2 => n6085, B1 => n5021, B2 => 
                           n6086, ZN => n6146);
   U6608 : AOI22_X1 port map( A1 => n204, A2 => n5022, B1 => n165, B2 => n5023,
                           ZN => n6144);
   U6609 : AOI22_X1 port map( A1 => n205, A2 => n5024, B1 => n162, B2 => n5025,
                           ZN => n6143);
   U6610 : NAND3_X1 port map( A1 => n6147, A2 => n6148, A3 => n6149, ZN => 
                           n12944);
   U6611 : AOI221_X1 port map( B1 => n151, B2 => n5029, C1 => n6083, C2 => 
                           MEM_IN(16), A => n6150, ZN => n6149);
   U6612 : OAI22_X1 port map( A1 => n11581, A2 => n6085, B1 => n5031, B2 => 
                           n6086, ZN => n6150);
   U6613 : AOI22_X1 port map( A1 => n204, A2 => n5032, B1 => n165, B2 => n5033,
                           ZN => n6148);
   U6614 : AOI22_X1 port map( A1 => n205, A2 => n5034, B1 => n162, B2 => n5035,
                           ZN => n6147);
   U6615 : NAND3_X1 port map( A1 => n6151, A2 => n6152, A3 => n6153, ZN => 
                           n12943);
   U6616 : AOI221_X1 port map( B1 => n151, B2 => n5039, C1 => n6083, C2 => 
                           MEM_IN(17), A => n6154, ZN => n6153);
   U6617 : OAI22_X1 port map( A1 => n11580, A2 => n6085, B1 => n5041, B2 => 
                           n6086, ZN => n6154);
   U6618 : AOI22_X1 port map( A1 => n204, A2 => n5042, B1 => n165, B2 => n5043,
                           ZN => n6152);
   U6619 : AOI22_X1 port map( A1 => n205, A2 => n5044, B1 => n162, B2 => n5045,
                           ZN => n6151);
   U6620 : NAND3_X1 port map( A1 => n6155, A2 => n6156, A3 => n6157, ZN => 
                           n12942);
   U6621 : AOI221_X1 port map( B1 => n151, B2 => n5049, C1 => n6083, C2 => 
                           MEM_IN(18), A => n6158, ZN => n6157);
   U6622 : OAI22_X1 port map( A1 => n11579, A2 => n6085, B1 => n5051, B2 => 
                           n6086, ZN => n6158);
   U6623 : AOI22_X1 port map( A1 => n204, A2 => n5052, B1 => n165, B2 => n5053,
                           ZN => n6156);
   U6624 : AOI22_X1 port map( A1 => n205, A2 => n5054, B1 => n162, B2 => n5055,
                           ZN => n6155);
   U6625 : NAND3_X1 port map( A1 => n6159, A2 => n6160, A3 => n6161, ZN => 
                           n12941);
   U6626 : AOI221_X1 port map( B1 => n151, B2 => n5059, C1 => n6083, C2 => 
                           MEM_IN(19), A => n6162, ZN => n6161);
   U6627 : OAI22_X1 port map( A1 => n11578, A2 => n6085, B1 => n5061, B2 => 
                           n6086, ZN => n6162);
   U6628 : AOI22_X1 port map( A1 => n204, A2 => n5062, B1 => n165, B2 => n5063,
                           ZN => n6160);
   U6629 : AOI22_X1 port map( A1 => n205, A2 => n5064, B1 => n162, B2 => n5065,
                           ZN => n6159);
   U6630 : NAND3_X1 port map( A1 => n6163, A2 => n6164, A3 => n6165, ZN => 
                           n12940);
   U6631 : AOI221_X1 port map( B1 => n151, B2 => n5069, C1 => n6083, C2 => 
                           MEM_IN(20), A => n6166, ZN => n6165);
   U6632 : OAI22_X1 port map( A1 => n11577, A2 => n6085, B1 => n5071, B2 => 
                           n6086, ZN => n6166);
   U6633 : AOI22_X1 port map( A1 => n204, A2 => n5072, B1 => n165, B2 => n5073,
                           ZN => n6164);
   U6634 : AOI22_X1 port map( A1 => n205, A2 => n5074, B1 => n162, B2 => n5075,
                           ZN => n6163);
   U6635 : NAND3_X1 port map( A1 => n6167, A2 => n6168, A3 => n6169, ZN => 
                           n12939);
   U6636 : AOI221_X1 port map( B1 => n151, B2 => n5079, C1 => n6083, C2 => 
                           MEM_IN(21), A => n6170, ZN => n6169);
   U6637 : OAI22_X1 port map( A1 => n11576, A2 => n6085, B1 => n5081, B2 => 
                           n6086, ZN => n6170);
   U6638 : AOI22_X1 port map( A1 => n204, A2 => n5082, B1 => n165, B2 => n5083,
                           ZN => n6168);
   U6639 : AOI22_X1 port map( A1 => n205, A2 => n5084, B1 => n162, B2 => n5085,
                           ZN => n6167);
   U6640 : NAND3_X1 port map( A1 => n6171, A2 => n6172, A3 => n6173, ZN => 
                           n12938);
   U6641 : AOI221_X1 port map( B1 => n151, B2 => n5089, C1 => n6083, C2 => 
                           MEM_IN(22), A => n6174, ZN => n6173);
   U6642 : OAI22_X1 port map( A1 => n11575, A2 => n6085, B1 => n5091, B2 => 
                           n6086, ZN => n6174);
   U6643 : AOI22_X1 port map( A1 => n204, A2 => n5092, B1 => n165, B2 => n5093,
                           ZN => n6172);
   U6644 : AOI22_X1 port map( A1 => n205, A2 => n5094, B1 => n162, B2 => n5095,
                           ZN => n6171);
   U6645 : NAND3_X1 port map( A1 => n6175, A2 => n6176, A3 => n6177, ZN => 
                           n12937);
   U6646 : AOI221_X1 port map( B1 => n151, B2 => n5099, C1 => n6083, C2 => 
                           MEM_IN(23), A => n6178, ZN => n6177);
   U6647 : OAI22_X1 port map( A1 => n11574, A2 => n6085, B1 => n5101, B2 => 
                           n6086, ZN => n6178);
   U6648 : AOI22_X1 port map( A1 => n204, A2 => n5102, B1 => n165, B2 => n5103,
                           ZN => n6176);
   U6649 : AOI22_X1 port map( A1 => n205, A2 => n5104, B1 => n162, B2 => n5105,
                           ZN => n6175);
   U6650 : NAND3_X1 port map( A1 => n6179, A2 => n6180, A3 => n6181, ZN => 
                           n12936);
   U6651 : AOI221_X1 port map( B1 => n151, B2 => n5109, C1 => n6083, C2 => 
                           MEM_IN(24), A => n6182, ZN => n6181);
   U6652 : OAI22_X1 port map( A1 => n11573, A2 => n6085, B1 => n5111, B2 => 
                           n6086, ZN => n6182);
   U6653 : AOI22_X1 port map( A1 => n204, A2 => n5112, B1 => n165, B2 => n5113,
                           ZN => n6180);
   U6654 : AOI22_X1 port map( A1 => n205, A2 => n5114, B1 => n162, B2 => n5115,
                           ZN => n6179);
   U6655 : NAND3_X1 port map( A1 => n6183, A2 => n6184, A3 => n6185, ZN => 
                           n12935);
   U6656 : AOI221_X1 port map( B1 => n151, B2 => n5119, C1 => n6083, C2 => 
                           MEM_IN(25), A => n6186, ZN => n6185);
   U6657 : OAI22_X1 port map( A1 => n11572, A2 => n6085, B1 => n5121, B2 => 
                           n6086, ZN => n6186);
   U6658 : AOI22_X1 port map( A1 => n204, A2 => n5122, B1 => n165, B2 => n5123,
                           ZN => n6184);
   U6659 : AOI22_X1 port map( A1 => n205, A2 => n5124, B1 => n162, B2 => n5125,
                           ZN => n6183);
   U6660 : NAND3_X1 port map( A1 => n6187, A2 => n6188, A3 => n6189, ZN => 
                           n12934);
   U6661 : AOI221_X1 port map( B1 => n151, B2 => n5129, C1 => n6083, C2 => 
                           MEM_IN(26), A => n6190, ZN => n6189);
   U6662 : OAI22_X1 port map( A1 => n11571, A2 => n6085, B1 => n5131, B2 => 
                           n6086, ZN => n6190);
   U6663 : AOI22_X1 port map( A1 => n204, A2 => n5132, B1 => n165, B2 => n5133,
                           ZN => n6188);
   U6664 : AOI22_X1 port map( A1 => n205, A2 => n5134, B1 => n162, B2 => n5135,
                           ZN => n6187);
   U6665 : NAND3_X1 port map( A1 => n6191, A2 => n6192, A3 => n6193, ZN => 
                           n12933);
   U6666 : AOI221_X1 port map( B1 => n151, B2 => n5139, C1 => n6083, C2 => 
                           MEM_IN(27), A => n6194, ZN => n6193);
   U6667 : OAI22_X1 port map( A1 => n11570, A2 => n6085, B1 => n5141, B2 => 
                           n6086, ZN => n6194);
   U6668 : AOI22_X1 port map( A1 => n204, A2 => n5142, B1 => n165, B2 => n5143,
                           ZN => n6192);
   U6669 : AOI22_X1 port map( A1 => n205, A2 => n5144, B1 => n162, B2 => n5145,
                           ZN => n6191);
   U6670 : NAND3_X1 port map( A1 => n6195, A2 => n6196, A3 => n6197, ZN => 
                           n12932);
   U6671 : AOI221_X1 port map( B1 => n151, B2 => n5149, C1 => n6083, C2 => 
                           MEM_IN(28), A => n6198, ZN => n6197);
   U6672 : OAI22_X1 port map( A1 => n11569, A2 => n6085, B1 => n5151, B2 => 
                           n6086, ZN => n6198);
   U6673 : AOI22_X1 port map( A1 => n204, A2 => n5152, B1 => n165, B2 => n5153,
                           ZN => n6196);
   U6674 : AOI22_X1 port map( A1 => n205, A2 => n5154, B1 => n162, B2 => n5155,
                           ZN => n6195);
   U6675 : NAND3_X1 port map( A1 => n6199, A2 => n6200, A3 => n6201, ZN => 
                           n12931);
   U6676 : AOI221_X1 port map( B1 => n151, B2 => n5159, C1 => n6083, C2 => 
                           MEM_IN(29), A => n6202, ZN => n6201);
   U6677 : OAI22_X1 port map( A1 => n11568, A2 => n6085, B1 => n5161, B2 => 
                           n6086, ZN => n6202);
   U6678 : AOI22_X1 port map( A1 => n204, A2 => n5162, B1 => n165, B2 => n5163,
                           ZN => n6200);
   U6679 : AOI22_X1 port map( A1 => n205, A2 => n5164, B1 => n162, B2 => n5165,
                           ZN => n6199);
   U6680 : NAND3_X1 port map( A1 => n6203, A2 => n6204, A3 => n6205, ZN => 
                           n12930);
   U6681 : AOI221_X1 port map( B1 => n151, B2 => n5169, C1 => n6083, C2 => 
                           MEM_IN(30), A => n6206, ZN => n6205);
   U6682 : OAI22_X1 port map( A1 => n11567, A2 => n6085, B1 => n5171, B2 => 
                           n6086, ZN => n6206);
   U6683 : AOI22_X1 port map( A1 => n204, A2 => n5172, B1 => n165, B2 => n5173,
                           ZN => n6204);
   U6684 : AOI22_X1 port map( A1 => n205, A2 => n5174, B1 => n162, B2 => n5175,
                           ZN => n6203);
   U6685 : NAND3_X1 port map( A1 => n6207, A2 => n6208, A3 => n6209, ZN => 
                           n12929);
   U6686 : AOI221_X1 port map( B1 => n151, B2 => n5179, C1 => n6083, C2 => 
                           MEM_IN(31), A => n6210, ZN => n6209);
   U6687 : OAI22_X1 port map( A1 => n11566, A2 => n6085, B1 => n5181, B2 => 
                           n6086, ZN => n6210);
   U6688 : AOI22_X1 port map( A1 => n204, A2 => n5191, B1 => n165, B2 => n5192,
                           ZN => n6208);
   U6689 : AOI22_X1 port map( A1 => n205, A2 => n5195, B1 => n162, B2 => n5196,
                           ZN => n6207);
   U6690 : AOI22_X1 port map( A1 => n6218, A2 => n6212, B1 => n4841, B2 => 
                           n6085, ZN => n6215);
   U6691 : NOR3_X1 port map( A1 => n4841, A2 => n6219, A3 => n6211, ZN => n6212
                           );
   U6692 : INV_X1 port map( A => n6085, ZN => n6219);
   U6693 : NOR2_X1 port map( A1 => n6211, A2 => n6213, ZN => n6221);
   U6694 : NAND2_X1 port map( A1 => n5767, A2 => n6222, ZN => n6211);
   U6695 : AOI211_X1 port map( C1 => n6223, C2 => n5208, A => n6214, B => RESET
                           , ZN => n6220);
   U6696 : OAI21_X1 port map( B1 => n5767, B2 => n4787, A => n6216, ZN => n6214
                           );
   U6697 : INV_X1 port map( A => n6224, ZN => n6216);
   U6698 : NOR3_X1 port map( A1 => n5371, A2 => n5525, A3 => n5214, ZN => n5767
                           );
   U6699 : INV_X1 port map( A => n6068, ZN => n5214);
   U6700 : INV_X1 port map( A => n6225, ZN => n5525);
   U6701 : INV_X1 port map( A => n5521, ZN => n5371);
   U6702 : INV_X1 port map( A => n6213, ZN => n6218);
   U6703 : NAND2_X1 port map( A1 => n6226, A2 => n6227, ZN => n6213);
   U6704 : INV_X1 port map( A => n5769, ZN => n5755);
   U6705 : NOR2_X1 port map( A1 => n6068, A2 => n4787, ZN => n5769);
   U6706 : NAND2_X1 port map( A1 => n6228, A2 => n5216, ZN => n6068);
   U6707 : NAND3_X1 port map( A1 => n6229, A2 => n6230, A3 => n6231, ZN => 
                           n12928);
   U6708 : AOI221_X1 port map( B1 => n6232, B2 => n4863, C1 => n6233, C2 => 
                           MEM_IN(0), A => n6234, ZN => n6231);
   U6709 : OAI22_X1 port map( A1 => n11565, A2 => n224, B1 => n4867, B2 => 
                           n6236, ZN => n6234);
   U6710 : AOI22_X1 port map( A1 => n6237, A2 => n4869, B1 => n6238, B2 => 
                           n4871, ZN => n6230);
   U6711 : AOI22_X1 port map( A1 => n6239, A2 => n4873, B1 => n6240, B2 => 
                           n4875, ZN => n6229);
   U6712 : NAND3_X1 port map( A1 => n6241, A2 => n6242, A3 => n6243, ZN => 
                           n12927);
   U6713 : AOI221_X1 port map( B1 => n6232, B2 => n4879, C1 => n6233, C2 => 
                           MEM_IN(1), A => n6244, ZN => n6243);
   U6714 : OAI22_X1 port map( A1 => n11564, A2 => n224, B1 => n4881, B2 => 
                           n6236, ZN => n6244);
   U6715 : AOI22_X1 port map( A1 => n6237, A2 => n4882, B1 => n6238, B2 => 
                           n4883, ZN => n6242);
   U6716 : AOI22_X1 port map( A1 => n6239, A2 => n4884, B1 => n6240, B2 => 
                           n4885, ZN => n6241);
   U6717 : NAND3_X1 port map( A1 => n6245, A2 => n6246, A3 => n6247, ZN => 
                           n12926);
   U6718 : AOI221_X1 port map( B1 => n6232, B2 => n4889, C1 => n6233, C2 => 
                           MEM_IN(2), A => n6248, ZN => n6247);
   U6719 : OAI22_X1 port map( A1 => n11563, A2 => n224, B1 => n4891, B2 => 
                           n6236, ZN => n6248);
   U6720 : AOI22_X1 port map( A1 => n6237, A2 => n4892, B1 => n6238, B2 => 
                           n4893, ZN => n6246);
   U6721 : AOI22_X1 port map( A1 => n6239, A2 => n4894, B1 => n6240, B2 => 
                           n4895, ZN => n6245);
   U6722 : NAND3_X1 port map( A1 => n6249, A2 => n6250, A3 => n6251, ZN => 
                           n12925);
   U6723 : AOI221_X1 port map( B1 => n6232, B2 => n4899, C1 => n6233, C2 => 
                           MEM_IN(3), A => n6252, ZN => n6251);
   U6724 : OAI22_X1 port map( A1 => n11562, A2 => n224, B1 => n4901, B2 => 
                           n6236, ZN => n6252);
   U6725 : AOI22_X1 port map( A1 => n6237, A2 => n4902, B1 => n6238, B2 => 
                           n4903, ZN => n6250);
   U6726 : AOI22_X1 port map( A1 => n6239, A2 => n4904, B1 => n6240, B2 => 
                           n4905, ZN => n6249);
   U6727 : NAND3_X1 port map( A1 => n6253, A2 => n6254, A3 => n6255, ZN => 
                           n12924);
   U6728 : AOI221_X1 port map( B1 => n6232, B2 => n4909, C1 => n6233, C2 => 
                           MEM_IN(4), A => n6256, ZN => n6255);
   U6729 : OAI22_X1 port map( A1 => n11561, A2 => n224, B1 => n4911, B2 => 
                           n6236, ZN => n6256);
   U6730 : AOI22_X1 port map( A1 => n6237, A2 => n4912, B1 => n6238, B2 => 
                           n4913, ZN => n6254);
   U6731 : AOI22_X1 port map( A1 => n6239, A2 => n4914, B1 => n6240, B2 => 
                           n4915, ZN => n6253);
   U6732 : NAND3_X1 port map( A1 => n6257, A2 => n6258, A3 => n6259, ZN => 
                           n12923);
   U6733 : AOI221_X1 port map( B1 => n6232, B2 => n4919, C1 => n6233, C2 => 
                           MEM_IN(5), A => n6260, ZN => n6259);
   U6734 : OAI22_X1 port map( A1 => n11560, A2 => n224, B1 => n4921, B2 => 
                           n6236, ZN => n6260);
   U6735 : AOI22_X1 port map( A1 => n6237, A2 => n4922, B1 => n6238, B2 => 
                           n4923, ZN => n6258);
   U6736 : AOI22_X1 port map( A1 => n6239, A2 => n4924, B1 => n6240, B2 => 
                           n4925, ZN => n6257);
   U6737 : NAND3_X1 port map( A1 => n6261, A2 => n6262, A3 => n6263, ZN => 
                           n12922);
   U6738 : AOI221_X1 port map( B1 => n6232, B2 => n4929, C1 => n6233, C2 => 
                           MEM_IN(6), A => n6264, ZN => n6263);
   U6739 : OAI22_X1 port map( A1 => n11559, A2 => n224, B1 => n4931, B2 => 
                           n6236, ZN => n6264);
   U6740 : AOI22_X1 port map( A1 => n6237, A2 => n4932, B1 => n6238, B2 => 
                           n4933, ZN => n6262);
   U6741 : AOI22_X1 port map( A1 => n6239, A2 => n4934, B1 => n6240, B2 => 
                           n4935, ZN => n6261);
   U6742 : NAND3_X1 port map( A1 => n6265, A2 => n6266, A3 => n6267, ZN => 
                           n12921);
   U6743 : AOI221_X1 port map( B1 => n6232, B2 => n4939, C1 => n6233, C2 => 
                           MEM_IN(7), A => n6268, ZN => n6267);
   U6744 : OAI22_X1 port map( A1 => n11558, A2 => n224, B1 => n4941, B2 => 
                           n6236, ZN => n6268);
   U6745 : AOI22_X1 port map( A1 => n6237, A2 => n4942, B1 => n6238, B2 => 
                           n4943, ZN => n6266);
   U6746 : AOI22_X1 port map( A1 => n6239, A2 => n4944, B1 => n6240, B2 => 
                           n4945, ZN => n6265);
   U6747 : NAND3_X1 port map( A1 => n6269, A2 => n6270, A3 => n6271, ZN => 
                           n12920);
   U6748 : AOI221_X1 port map( B1 => n6232, B2 => n4949, C1 => n6233, C2 => 
                           MEM_IN(8), A => n6272, ZN => n6271);
   U6749 : OAI22_X1 port map( A1 => n11557, A2 => n224, B1 => n4951, B2 => 
                           n6236, ZN => n6272);
   U6750 : AOI22_X1 port map( A1 => n6237, A2 => n4952, B1 => n6238, B2 => 
                           n4953, ZN => n6270);
   U6751 : AOI22_X1 port map( A1 => n6239, A2 => n4954, B1 => n6240, B2 => 
                           n4955, ZN => n6269);
   U6752 : NAND3_X1 port map( A1 => n6273, A2 => n6274, A3 => n6275, ZN => 
                           n12919);
   U6753 : AOI221_X1 port map( B1 => n6232, B2 => n4959, C1 => n6233, C2 => 
                           MEM_IN(9), A => n6276, ZN => n6275);
   U6754 : OAI22_X1 port map( A1 => n11556, A2 => n224, B1 => n4961, B2 => 
                           n6236, ZN => n6276);
   U6755 : AOI22_X1 port map( A1 => n6237, A2 => n4962, B1 => n6238, B2 => 
                           n4963, ZN => n6274);
   U6756 : AOI22_X1 port map( A1 => n6239, A2 => n4964, B1 => n6240, B2 => 
                           n4965, ZN => n6273);
   U6757 : NAND3_X1 port map( A1 => n6277, A2 => n6278, A3 => n6279, ZN => 
                           n12918);
   U6758 : AOI221_X1 port map( B1 => n6232, B2 => n4969, C1 => n6233, C2 => 
                           MEM_IN(10), A => n6280, ZN => n6279);
   U6759 : OAI22_X1 port map( A1 => n11555, A2 => n224, B1 => n4971, B2 => 
                           n6236, ZN => n6280);
   U6760 : AOI22_X1 port map( A1 => n6237, A2 => n4972, B1 => n6238, B2 => 
                           n4973, ZN => n6278);
   U6761 : AOI22_X1 port map( A1 => n6239, A2 => n4974, B1 => n6240, B2 => 
                           n4975, ZN => n6277);
   U6762 : NAND3_X1 port map( A1 => n6281, A2 => n6282, A3 => n6283, ZN => 
                           n12917);
   U6763 : AOI221_X1 port map( B1 => n6232, B2 => n4979, C1 => n6233, C2 => 
                           MEM_IN(11), A => n6284, ZN => n6283);
   U6764 : OAI22_X1 port map( A1 => n11554, A2 => n224, B1 => n4981, B2 => 
                           n6236, ZN => n6284);
   U6765 : AOI22_X1 port map( A1 => n6237, A2 => n4982, B1 => n6238, B2 => 
                           n4983, ZN => n6282);
   U6766 : AOI22_X1 port map( A1 => n6239, A2 => n4984, B1 => n6240, B2 => 
                           n4985, ZN => n6281);
   U6767 : NAND3_X1 port map( A1 => n6285, A2 => n6286, A3 => n6287, ZN => 
                           n12916);
   U6768 : AOI221_X1 port map( B1 => n6232, B2 => n4989, C1 => n6233, C2 => 
                           MEM_IN(12), A => n6288, ZN => n6287);
   U6769 : OAI22_X1 port map( A1 => n11553, A2 => n224, B1 => n4991, B2 => 
                           n6236, ZN => n6288);
   U6770 : AOI22_X1 port map( A1 => n6237, A2 => n4992, B1 => n6238, B2 => 
                           n4993, ZN => n6286);
   U6771 : AOI22_X1 port map( A1 => n6239, A2 => n4994, B1 => n6240, B2 => 
                           n4995, ZN => n6285);
   U6772 : NAND3_X1 port map( A1 => n6289, A2 => n6290, A3 => n6291, ZN => 
                           n12915);
   U6773 : AOI221_X1 port map( B1 => n6232, B2 => n4999, C1 => n6233, C2 => 
                           MEM_IN(13), A => n6292, ZN => n6291);
   U6774 : OAI22_X1 port map( A1 => n11552, A2 => n224, B1 => n5001, B2 => 
                           n6236, ZN => n6292);
   U6775 : AOI22_X1 port map( A1 => n6237, A2 => n5002, B1 => n6238, B2 => 
                           n5003, ZN => n6290);
   U6776 : AOI22_X1 port map( A1 => n6239, A2 => n5004, B1 => n6240, B2 => 
                           n5005, ZN => n6289);
   U6777 : NAND3_X1 port map( A1 => n6293, A2 => n6294, A3 => n6295, ZN => 
                           n12914);
   U6778 : AOI221_X1 port map( B1 => n6232, B2 => n5009, C1 => n6233, C2 => 
                           MEM_IN(14), A => n6296, ZN => n6295);
   U6779 : OAI22_X1 port map( A1 => n11551, A2 => n224, B1 => n5011, B2 => 
                           n6236, ZN => n6296);
   U6780 : AOI22_X1 port map( A1 => n6237, A2 => n5012, B1 => n6238, B2 => 
                           n5013, ZN => n6294);
   U6781 : AOI22_X1 port map( A1 => n6239, A2 => n5014, B1 => n6240, B2 => 
                           n5015, ZN => n6293);
   U6782 : NAND3_X1 port map( A1 => n6297, A2 => n6298, A3 => n6299, ZN => 
                           n12913);
   U6783 : AOI221_X1 port map( B1 => n6232, B2 => n5019, C1 => n6233, C2 => 
                           MEM_IN(15), A => n6300, ZN => n6299);
   U6784 : OAI22_X1 port map( A1 => n11550, A2 => n224, B1 => n5021, B2 => 
                           n6236, ZN => n6300);
   U6785 : AOI22_X1 port map( A1 => n6237, A2 => n5022, B1 => n6238, B2 => 
                           n5023, ZN => n6298);
   U6786 : AOI22_X1 port map( A1 => n6239, A2 => n5024, B1 => n6240, B2 => 
                           n5025, ZN => n6297);
   U6787 : NAND3_X1 port map( A1 => n6301, A2 => n6302, A3 => n6303, ZN => 
                           n12912);
   U6788 : AOI221_X1 port map( B1 => n6232, B2 => n5029, C1 => n6233, C2 => 
                           MEM_IN(16), A => n6304, ZN => n6303);
   U6789 : OAI22_X1 port map( A1 => n11549, A2 => n224, B1 => n5031, B2 => 
                           n6236, ZN => n6304);
   U6790 : AOI22_X1 port map( A1 => n6237, A2 => n5032, B1 => n6238, B2 => 
                           n5033, ZN => n6302);
   U6791 : AOI22_X1 port map( A1 => n6239, A2 => n5034, B1 => n6240, B2 => 
                           n5035, ZN => n6301);
   U6792 : NAND3_X1 port map( A1 => n6305, A2 => n6306, A3 => n6307, ZN => 
                           n12911);
   U6793 : AOI221_X1 port map( B1 => n6232, B2 => n5039, C1 => n6233, C2 => 
                           MEM_IN(17), A => n6308, ZN => n6307);
   U6794 : OAI22_X1 port map( A1 => n11548, A2 => n224, B1 => n5041, B2 => 
                           n6236, ZN => n6308);
   U6795 : AOI22_X1 port map( A1 => n6237, A2 => n5042, B1 => n6238, B2 => 
                           n5043, ZN => n6306);
   U6796 : AOI22_X1 port map( A1 => n6239, A2 => n5044, B1 => n6240, B2 => 
                           n5045, ZN => n6305);
   U6797 : NAND3_X1 port map( A1 => n6309, A2 => n6310, A3 => n6311, ZN => 
                           n12910);
   U6798 : AOI221_X1 port map( B1 => n6232, B2 => n5049, C1 => n6233, C2 => 
                           MEM_IN(18), A => n6312, ZN => n6311);
   U6799 : OAI22_X1 port map( A1 => n11547, A2 => n224, B1 => n5051, B2 => 
                           n6236, ZN => n6312);
   U6800 : AOI22_X1 port map( A1 => n6237, A2 => n5052, B1 => n6238, B2 => 
                           n5053, ZN => n6310);
   U6801 : AOI22_X1 port map( A1 => n6239, A2 => n5054, B1 => n6240, B2 => 
                           n5055, ZN => n6309);
   U6802 : NAND3_X1 port map( A1 => n6313, A2 => n6314, A3 => n6315, ZN => 
                           n12909);
   U6803 : AOI221_X1 port map( B1 => n6232, B2 => n5059, C1 => n6233, C2 => 
                           MEM_IN(19), A => n6316, ZN => n6315);
   U6804 : OAI22_X1 port map( A1 => n11546, A2 => n224, B1 => n5061, B2 => 
                           n6236, ZN => n6316);
   U6805 : AOI22_X1 port map( A1 => n6237, A2 => n5062, B1 => n6238, B2 => 
                           n5063, ZN => n6314);
   U6806 : AOI22_X1 port map( A1 => n6239, A2 => n5064, B1 => n6240, B2 => 
                           n5065, ZN => n6313);
   U6807 : NAND3_X1 port map( A1 => n6317, A2 => n6318, A3 => n6319, ZN => 
                           n12908);
   U6808 : AOI221_X1 port map( B1 => n6232, B2 => n5069, C1 => n6233, C2 => 
                           MEM_IN(20), A => n6320, ZN => n6319);
   U6809 : OAI22_X1 port map( A1 => n11545, A2 => n224, B1 => n5071, B2 => 
                           n6236, ZN => n6320);
   U6810 : AOI22_X1 port map( A1 => n6237, A2 => n5072, B1 => n6238, B2 => 
                           n5073, ZN => n6318);
   U6811 : AOI22_X1 port map( A1 => n6239, A2 => n5074, B1 => n6240, B2 => 
                           n5075, ZN => n6317);
   U6812 : NAND3_X1 port map( A1 => n6321, A2 => n6322, A3 => n6323, ZN => 
                           n12907);
   U6813 : AOI221_X1 port map( B1 => n6232, B2 => n5079, C1 => n6233, C2 => 
                           MEM_IN(21), A => n6324, ZN => n6323);
   U6814 : OAI22_X1 port map( A1 => n11544, A2 => n224, B1 => n5081, B2 => 
                           n6236, ZN => n6324);
   U6815 : AOI22_X1 port map( A1 => n6237, A2 => n5082, B1 => n6238, B2 => 
                           n5083, ZN => n6322);
   U6816 : AOI22_X1 port map( A1 => n6239, A2 => n5084, B1 => n6240, B2 => 
                           n5085, ZN => n6321);
   U6817 : NAND3_X1 port map( A1 => n6325, A2 => n6326, A3 => n6327, ZN => 
                           n12906);
   U6818 : AOI221_X1 port map( B1 => n6232, B2 => n5089, C1 => n6233, C2 => 
                           MEM_IN(22), A => n6328, ZN => n6327);
   U6819 : OAI22_X1 port map( A1 => n11543, A2 => n224, B1 => n5091, B2 => 
                           n6236, ZN => n6328);
   U6820 : AOI22_X1 port map( A1 => n6237, A2 => n5092, B1 => n6238, B2 => 
                           n5093, ZN => n6326);
   U6821 : AOI22_X1 port map( A1 => n6239, A2 => n5094, B1 => n6240, B2 => 
                           n5095, ZN => n6325);
   U6822 : NAND3_X1 port map( A1 => n6329, A2 => n6330, A3 => n6331, ZN => 
                           n12905);
   U6823 : AOI221_X1 port map( B1 => n6232, B2 => n5099, C1 => n6233, C2 => 
                           MEM_IN(23), A => n6332, ZN => n6331);
   U6824 : OAI22_X1 port map( A1 => n11542, A2 => n224, B1 => n5101, B2 => 
                           n6236, ZN => n6332);
   U6825 : AOI22_X1 port map( A1 => n6237, A2 => n5102, B1 => n6238, B2 => 
                           n5103, ZN => n6330);
   U6826 : AOI22_X1 port map( A1 => n6239, A2 => n5104, B1 => n6240, B2 => 
                           n5105, ZN => n6329);
   U6827 : NAND3_X1 port map( A1 => n6333, A2 => n6334, A3 => n6335, ZN => 
                           n12904);
   U6828 : AOI221_X1 port map( B1 => n6232, B2 => n5109, C1 => n6233, C2 => 
                           MEM_IN(24), A => n6336, ZN => n6335);
   U6829 : OAI22_X1 port map( A1 => n11541, A2 => n224, B1 => n5111, B2 => 
                           n6236, ZN => n6336);
   U6830 : AOI22_X1 port map( A1 => n6237, A2 => n5112, B1 => n6238, B2 => 
                           n5113, ZN => n6334);
   U6831 : AOI22_X1 port map( A1 => n6239, A2 => n5114, B1 => n6240, B2 => 
                           n5115, ZN => n6333);
   U6832 : NAND3_X1 port map( A1 => n6337, A2 => n6338, A3 => n6339, ZN => 
                           n12903);
   U6833 : AOI221_X1 port map( B1 => n6232, B2 => n5119, C1 => n6233, C2 => 
                           MEM_IN(25), A => n6340, ZN => n6339);
   U6834 : OAI22_X1 port map( A1 => n11540, A2 => n224, B1 => n5121, B2 => 
                           n6236, ZN => n6340);
   U6835 : AOI22_X1 port map( A1 => n6237, A2 => n5122, B1 => n6238, B2 => 
                           n5123, ZN => n6338);
   U6836 : AOI22_X1 port map( A1 => n6239, A2 => n5124, B1 => n6240, B2 => 
                           n5125, ZN => n6337);
   U6837 : NAND3_X1 port map( A1 => n6341, A2 => n6342, A3 => n6343, ZN => 
                           n12902);
   U6838 : AOI221_X1 port map( B1 => n6232, B2 => n5129, C1 => n6233, C2 => 
                           MEM_IN(26), A => n6344, ZN => n6343);
   U6839 : OAI22_X1 port map( A1 => n11539, A2 => n224, B1 => n5131, B2 => 
                           n6236, ZN => n6344);
   U6840 : AOI22_X1 port map( A1 => n6237, A2 => n5132, B1 => n6238, B2 => 
                           n5133, ZN => n6342);
   U6841 : AOI22_X1 port map( A1 => n6239, A2 => n5134, B1 => n6240, B2 => 
                           n5135, ZN => n6341);
   U6842 : NAND3_X1 port map( A1 => n6345, A2 => n6346, A3 => n6347, ZN => 
                           n12901);
   U6843 : AOI221_X1 port map( B1 => n6232, B2 => n5139, C1 => n6233, C2 => 
                           MEM_IN(27), A => n6348, ZN => n6347);
   U6844 : OAI22_X1 port map( A1 => n11538, A2 => n224, B1 => n5141, B2 => 
                           n6236, ZN => n6348);
   U6845 : AOI22_X1 port map( A1 => n6237, A2 => n5142, B1 => n6238, B2 => 
                           n5143, ZN => n6346);
   U6846 : AOI22_X1 port map( A1 => n6239, A2 => n5144, B1 => n6240, B2 => 
                           n5145, ZN => n6345);
   U6847 : NAND3_X1 port map( A1 => n6349, A2 => n6350, A3 => n6351, ZN => 
                           n12900);
   U6848 : AOI221_X1 port map( B1 => n6232, B2 => n5149, C1 => n6233, C2 => 
                           MEM_IN(28), A => n6352, ZN => n6351);
   U6849 : OAI22_X1 port map( A1 => n11537, A2 => n224, B1 => n5151, B2 => 
                           n6236, ZN => n6352);
   U6850 : AOI22_X1 port map( A1 => n6237, A2 => n5152, B1 => n6238, B2 => 
                           n5153, ZN => n6350);
   U6851 : AOI22_X1 port map( A1 => n6239, A2 => n5154, B1 => n6240, B2 => 
                           n5155, ZN => n6349);
   U6852 : NAND3_X1 port map( A1 => n6353, A2 => n6354, A3 => n6355, ZN => 
                           n12899);
   U6853 : AOI221_X1 port map( B1 => n6232, B2 => n5159, C1 => n6233, C2 => 
                           MEM_IN(29), A => n6356, ZN => n6355);
   U6854 : OAI22_X1 port map( A1 => n11536, A2 => n224, B1 => n5161, B2 => 
                           n6236, ZN => n6356);
   U6855 : AOI22_X1 port map( A1 => n6237, A2 => n5162, B1 => n6238, B2 => 
                           n5163, ZN => n6354);
   U6856 : AOI22_X1 port map( A1 => n6239, A2 => n5164, B1 => n6240, B2 => 
                           n5165, ZN => n6353);
   U6857 : NAND3_X1 port map( A1 => n6357, A2 => n6358, A3 => n6359, ZN => 
                           n12898);
   U6858 : AOI221_X1 port map( B1 => n6232, B2 => n5169, C1 => n6233, C2 => 
                           MEM_IN(30), A => n6360, ZN => n6359);
   U6859 : OAI22_X1 port map( A1 => n11535, A2 => n224, B1 => n5171, B2 => 
                           n6236, ZN => n6360);
   U6860 : AOI22_X1 port map( A1 => n6237, A2 => n5172, B1 => n6238, B2 => 
                           n5173, ZN => n6358);
   U6861 : AOI22_X1 port map( A1 => n6239, A2 => n5174, B1 => n6240, B2 => 
                           n5175, ZN => n6357);
   U6862 : NAND3_X1 port map( A1 => n6361, A2 => n6362, A3 => n6363, ZN => 
                           n12897);
   U6863 : AOI221_X1 port map( B1 => n6232, B2 => n5179, C1 => n6233, C2 => 
                           MEM_IN(31), A => n6364, ZN => n6363);
   U6864 : OAI22_X1 port map( A1 => n11534, A2 => n224, B1 => n5181, B2 => 
                           n6236, ZN => n6364);
   U6865 : AOI22_X1 port map( A1 => n6237, A2 => n5191, B1 => n6238, B2 => 
                           n5192, ZN => n6362);
   U6866 : AOI22_X1 port map( A1 => n6239, A2 => n5195, B1 => n6240, B2 => 
                           n5196, ZN => n6361);
   U6867 : OAI22_X1 port map( A1 => n6366, A2 => n6370, B1 => n208, B2 => n223,
                           ZN => n6367);
   U6868 : INV_X1 port map( A => n6365, ZN => n6370);
   U6869 : NOR3_X1 port map( A1 => n5213, A2 => n223, A3 => n4841, ZN => n6365)
                           ;
   U6870 : OAI22_X1 port map( A1 => n4786, A2 => n6371, B1 => n6372, B2 => 
                           n5204, ZN => n6235);
   U6871 : NOR2_X1 port map( A1 => n5213, A2 => n6366, ZN => n6372);
   U6872 : NOR4_X1 port map( A1 => n6373, A2 => n6224, A3 => RESET, A4 => n6369
                           , ZN => n6371);
   U6873 : OAI211_X1 port map( C1 => n5770, C2 => n6374, A => n6217, B => n6066
                           , ZN => n6373);
   U6874 : INV_X1 port map( A => n5917, ZN => n6217);
   U6875 : INV_X1 port map( A => n5208, ZN => n5770);
   U6876 : NOR4_X1 port map( A1 => n6375, A2 => n6376, A3 => n6377, A4 => n6378
                           , ZN => n5208);
   U6877 : INV_X1 port map( A => WR, ZN => n6375);
   U6878 : NAND4_X1 port map( A1 => n6222, A2 => n5521, A3 => n6225, A4 => 
                           n6227, ZN => n5213);
   U6879 : NAND2_X1 port map( A1 => n6379, A2 => n6380, ZN => n6366);
   U6880 : NOR2_X1 port map( A1 => n5521, A2 => n4787, ZN => n5917);
   U6881 : NAND2_X1 port map( A1 => n6381, A2 => n5216, ZN => n5521);
   U6882 : NAND3_X1 port map( A1 => n6382, A2 => n6383, A3 => n6384, ZN => 
                           n12896);
   U6883 : AOI221_X1 port map( B1 => n6385, B2 => n4863, C1 => n6386, C2 => 
                           MEM_IN(0), A => n6387, ZN => n6384);
   U6884 : OAI22_X1 port map( A1 => n11533, A2 => n226, B1 => n4867, B2 => 
                           n6389, ZN => n6387);
   U6885 : AOI22_X1 port map( A1 => n6390, A2 => n4869, B1 => n6391, B2 => 
                           n4871, ZN => n6383);
   U6886 : AOI22_X1 port map( A1 => n6392, A2 => n4873, B1 => n6393, B2 => 
                           n4875, ZN => n6382);
   U6887 : NAND3_X1 port map( A1 => n6394, A2 => n6395, A3 => n6396, ZN => 
                           n12895);
   U6888 : AOI221_X1 port map( B1 => n6385, B2 => n4879, C1 => n6386, C2 => 
                           MEM_IN(1), A => n6397, ZN => n6396);
   U6889 : OAI22_X1 port map( A1 => n11532, A2 => n226, B1 => n4881, B2 => 
                           n6389, ZN => n6397);
   U6890 : AOI22_X1 port map( A1 => n6390, A2 => n4882, B1 => n6391, B2 => 
                           n4883, ZN => n6395);
   U6891 : AOI22_X1 port map( A1 => n6392, A2 => n4884, B1 => n6393, B2 => 
                           n4885, ZN => n6394);
   U6892 : NAND3_X1 port map( A1 => n6398, A2 => n6399, A3 => n6400, ZN => 
                           n12894);
   U6893 : AOI221_X1 port map( B1 => n6385, B2 => n4889, C1 => n6386, C2 => 
                           MEM_IN(2), A => n6401, ZN => n6400);
   U6894 : OAI22_X1 port map( A1 => n11531, A2 => n226, B1 => n4891, B2 => 
                           n6389, ZN => n6401);
   U6895 : AOI22_X1 port map( A1 => n6390, A2 => n4892, B1 => n6391, B2 => 
                           n4893, ZN => n6399);
   U6896 : AOI22_X1 port map( A1 => n6392, A2 => n4894, B1 => n6393, B2 => 
                           n4895, ZN => n6398);
   U6897 : NAND3_X1 port map( A1 => n6402, A2 => n6403, A3 => n6404, ZN => 
                           n12893);
   U6898 : AOI221_X1 port map( B1 => n6385, B2 => n4899, C1 => n6386, C2 => 
                           MEM_IN(3), A => n6405, ZN => n6404);
   U6899 : OAI22_X1 port map( A1 => n11530, A2 => n226, B1 => n4901, B2 => 
                           n6389, ZN => n6405);
   U6900 : AOI22_X1 port map( A1 => n6390, A2 => n4902, B1 => n6391, B2 => 
                           n4903, ZN => n6403);
   U6901 : AOI22_X1 port map( A1 => n6392, A2 => n4904, B1 => n6393, B2 => 
                           n4905, ZN => n6402);
   U6902 : NAND3_X1 port map( A1 => n6406, A2 => n6407, A3 => n6408, ZN => 
                           n12892);
   U6903 : AOI221_X1 port map( B1 => n6385, B2 => n4909, C1 => n6386, C2 => 
                           MEM_IN(4), A => n6409, ZN => n6408);
   U6904 : OAI22_X1 port map( A1 => n11529, A2 => n226, B1 => n4911, B2 => 
                           n6389, ZN => n6409);
   U6905 : AOI22_X1 port map( A1 => n6390, A2 => n4912, B1 => n6391, B2 => 
                           n4913, ZN => n6407);
   U6906 : AOI22_X1 port map( A1 => n6392, A2 => n4914, B1 => n6393, B2 => 
                           n4915, ZN => n6406);
   U6907 : NAND3_X1 port map( A1 => n6410, A2 => n6411, A3 => n6412, ZN => 
                           n12891);
   U6908 : AOI221_X1 port map( B1 => n6385, B2 => n4919, C1 => n6386, C2 => 
                           MEM_IN(5), A => n6413, ZN => n6412);
   U6909 : OAI22_X1 port map( A1 => n11528, A2 => n226, B1 => n4921, B2 => 
                           n6389, ZN => n6413);
   U6910 : AOI22_X1 port map( A1 => n6390, A2 => n4922, B1 => n6391, B2 => 
                           n4923, ZN => n6411);
   U6911 : AOI22_X1 port map( A1 => n6392, A2 => n4924, B1 => n6393, B2 => 
                           n4925, ZN => n6410);
   U6912 : NAND3_X1 port map( A1 => n6414, A2 => n6415, A3 => n6416, ZN => 
                           n12890);
   U6913 : AOI221_X1 port map( B1 => n6385, B2 => n4929, C1 => n6386, C2 => 
                           MEM_IN(6), A => n6417, ZN => n6416);
   U6914 : OAI22_X1 port map( A1 => n11527, A2 => n226, B1 => n4931, B2 => 
                           n6389, ZN => n6417);
   U6915 : AOI22_X1 port map( A1 => n6390, A2 => n4932, B1 => n6391, B2 => 
                           n4933, ZN => n6415);
   U6916 : AOI22_X1 port map( A1 => n6392, A2 => n4934, B1 => n6393, B2 => 
                           n4935, ZN => n6414);
   U6917 : NAND3_X1 port map( A1 => n6418, A2 => n6419, A3 => n6420, ZN => 
                           n12889);
   U6918 : AOI221_X1 port map( B1 => n6385, B2 => n4939, C1 => n6386, C2 => 
                           MEM_IN(7), A => n6421, ZN => n6420);
   U6919 : OAI22_X1 port map( A1 => n11526, A2 => n226, B1 => n4941, B2 => 
                           n6389, ZN => n6421);
   U6920 : AOI22_X1 port map( A1 => n6390, A2 => n4942, B1 => n6391, B2 => 
                           n4943, ZN => n6419);
   U6921 : AOI22_X1 port map( A1 => n6392, A2 => n4944, B1 => n6393, B2 => 
                           n4945, ZN => n6418);
   U6922 : NAND3_X1 port map( A1 => n6422, A2 => n6423, A3 => n6424, ZN => 
                           n12888);
   U6923 : AOI221_X1 port map( B1 => n6385, B2 => n4949, C1 => n6386, C2 => 
                           MEM_IN(8), A => n6425, ZN => n6424);
   U6924 : OAI22_X1 port map( A1 => n11525, A2 => n226, B1 => n4951, B2 => 
                           n6389, ZN => n6425);
   U6925 : AOI22_X1 port map( A1 => n6390, A2 => n4952, B1 => n6391, B2 => 
                           n4953, ZN => n6423);
   U6926 : AOI22_X1 port map( A1 => n6392, A2 => n4954, B1 => n6393, B2 => 
                           n4955, ZN => n6422);
   U6927 : NAND3_X1 port map( A1 => n6426, A2 => n6427, A3 => n6428, ZN => 
                           n12887);
   U6928 : AOI221_X1 port map( B1 => n6385, B2 => n4959, C1 => n6386, C2 => 
                           MEM_IN(9), A => n6429, ZN => n6428);
   U6929 : OAI22_X1 port map( A1 => n11524, A2 => n226, B1 => n4961, B2 => 
                           n6389, ZN => n6429);
   U6930 : AOI22_X1 port map( A1 => n6390, A2 => n4962, B1 => n6391, B2 => 
                           n4963, ZN => n6427);
   U6931 : AOI22_X1 port map( A1 => n6392, A2 => n4964, B1 => n6393, B2 => 
                           n4965, ZN => n6426);
   U6932 : NAND3_X1 port map( A1 => n6430, A2 => n6431, A3 => n6432, ZN => 
                           n12886);
   U6933 : AOI221_X1 port map( B1 => n6385, B2 => n4969, C1 => n6386, C2 => 
                           MEM_IN(10), A => n6433, ZN => n6432);
   U6934 : OAI22_X1 port map( A1 => n11523, A2 => n226, B1 => n4971, B2 => 
                           n6389, ZN => n6433);
   U6935 : AOI22_X1 port map( A1 => n6390, A2 => n4972, B1 => n6391, B2 => 
                           n4973, ZN => n6431);
   U6936 : AOI22_X1 port map( A1 => n6392, A2 => n4974, B1 => n6393, B2 => 
                           n4975, ZN => n6430);
   U6937 : NAND3_X1 port map( A1 => n6434, A2 => n6435, A3 => n6436, ZN => 
                           n12885);
   U6938 : AOI221_X1 port map( B1 => n6385, B2 => n4979, C1 => n6386, C2 => 
                           MEM_IN(11), A => n6437, ZN => n6436);
   U6939 : OAI22_X1 port map( A1 => n11522, A2 => n226, B1 => n4981, B2 => 
                           n6389, ZN => n6437);
   U6940 : AOI22_X1 port map( A1 => n6390, A2 => n4982, B1 => n6391, B2 => 
                           n4983, ZN => n6435);
   U6941 : AOI22_X1 port map( A1 => n6392, A2 => n4984, B1 => n6393, B2 => 
                           n4985, ZN => n6434);
   U6942 : NAND3_X1 port map( A1 => n6438, A2 => n6439, A3 => n6440, ZN => 
                           n12884);
   U6943 : AOI221_X1 port map( B1 => n6385, B2 => n4989, C1 => n6386, C2 => 
                           MEM_IN(12), A => n6441, ZN => n6440);
   U6944 : OAI22_X1 port map( A1 => n11521, A2 => n226, B1 => n4991, B2 => 
                           n6389, ZN => n6441);
   U6945 : AOI22_X1 port map( A1 => n6390, A2 => n4992, B1 => n6391, B2 => 
                           n4993, ZN => n6439);
   U6946 : AOI22_X1 port map( A1 => n6392, A2 => n4994, B1 => n6393, B2 => 
                           n4995, ZN => n6438);
   U6947 : NAND3_X1 port map( A1 => n6442, A2 => n6443, A3 => n6444, ZN => 
                           n12883);
   U6948 : AOI221_X1 port map( B1 => n6385, B2 => n4999, C1 => n6386, C2 => 
                           MEM_IN(13), A => n6445, ZN => n6444);
   U6949 : OAI22_X1 port map( A1 => n11520, A2 => n226, B1 => n5001, B2 => 
                           n6389, ZN => n6445);
   U6950 : AOI22_X1 port map( A1 => n6390, A2 => n5002, B1 => n6391, B2 => 
                           n5003, ZN => n6443);
   U6951 : AOI22_X1 port map( A1 => n6392, A2 => n5004, B1 => n6393, B2 => 
                           n5005, ZN => n6442);
   U6952 : NAND3_X1 port map( A1 => n6446, A2 => n6447, A3 => n6448, ZN => 
                           n12882);
   U6953 : AOI221_X1 port map( B1 => n6385, B2 => n5009, C1 => n6386, C2 => 
                           MEM_IN(14), A => n6449, ZN => n6448);
   U6954 : OAI22_X1 port map( A1 => n11519, A2 => n226, B1 => n5011, B2 => 
                           n6389, ZN => n6449);
   U6955 : AOI22_X1 port map( A1 => n6390, A2 => n5012, B1 => n6391, B2 => 
                           n5013, ZN => n6447);
   U6956 : AOI22_X1 port map( A1 => n6392, A2 => n5014, B1 => n6393, B2 => 
                           n5015, ZN => n6446);
   U6957 : NAND3_X1 port map( A1 => n6450, A2 => n6451, A3 => n6452, ZN => 
                           n12881);
   U6958 : AOI221_X1 port map( B1 => n6385, B2 => n5019, C1 => n6386, C2 => 
                           MEM_IN(15), A => n6453, ZN => n6452);
   U6959 : OAI22_X1 port map( A1 => n11518, A2 => n226, B1 => n5021, B2 => 
                           n6389, ZN => n6453);
   U6960 : AOI22_X1 port map( A1 => n6390, A2 => n5022, B1 => n6391, B2 => 
                           n5023, ZN => n6451);
   U6961 : AOI22_X1 port map( A1 => n6392, A2 => n5024, B1 => n6393, B2 => 
                           n5025, ZN => n6450);
   U6962 : NAND3_X1 port map( A1 => n6454, A2 => n6455, A3 => n6456, ZN => 
                           n12880);
   U6963 : AOI221_X1 port map( B1 => n6385, B2 => n5029, C1 => n6386, C2 => 
                           MEM_IN(16), A => n6457, ZN => n6456);
   U6964 : OAI22_X1 port map( A1 => n11517, A2 => n226, B1 => n5031, B2 => 
                           n6389, ZN => n6457);
   U6965 : AOI22_X1 port map( A1 => n6390, A2 => n5032, B1 => n6391, B2 => 
                           n5033, ZN => n6455);
   U6966 : AOI22_X1 port map( A1 => n6392, A2 => n5034, B1 => n6393, B2 => 
                           n5035, ZN => n6454);
   U6967 : NAND3_X1 port map( A1 => n6458, A2 => n6459, A3 => n6460, ZN => 
                           n12879);
   U6968 : AOI221_X1 port map( B1 => n6385, B2 => n5039, C1 => n6386, C2 => 
                           MEM_IN(17), A => n6461, ZN => n6460);
   U6969 : OAI22_X1 port map( A1 => n11516, A2 => n226, B1 => n5041, B2 => 
                           n6389, ZN => n6461);
   U6970 : AOI22_X1 port map( A1 => n6390, A2 => n5042, B1 => n6391, B2 => 
                           n5043, ZN => n6459);
   U6971 : AOI22_X1 port map( A1 => n6392, A2 => n5044, B1 => n6393, B2 => 
                           n5045, ZN => n6458);
   U6972 : NAND3_X1 port map( A1 => n6462, A2 => n6463, A3 => n6464, ZN => 
                           n12878);
   U6973 : AOI221_X1 port map( B1 => n6385, B2 => n5049, C1 => n6386, C2 => 
                           MEM_IN(18), A => n6465, ZN => n6464);
   U6974 : OAI22_X1 port map( A1 => n11515, A2 => n226, B1 => n5051, B2 => 
                           n6389, ZN => n6465);
   U6975 : AOI22_X1 port map( A1 => n6390, A2 => n5052, B1 => n6391, B2 => 
                           n5053, ZN => n6463);
   U6976 : AOI22_X1 port map( A1 => n6392, A2 => n5054, B1 => n6393, B2 => 
                           n5055, ZN => n6462);
   U6977 : NAND3_X1 port map( A1 => n6466, A2 => n6467, A3 => n6468, ZN => 
                           n12877);
   U6978 : AOI221_X1 port map( B1 => n6385, B2 => n5059, C1 => n6386, C2 => 
                           MEM_IN(19), A => n6469, ZN => n6468);
   U6979 : OAI22_X1 port map( A1 => n11514, A2 => n226, B1 => n5061, B2 => 
                           n6389, ZN => n6469);
   U6980 : AOI22_X1 port map( A1 => n6390, A2 => n5062, B1 => n6391, B2 => 
                           n5063, ZN => n6467);
   U6981 : AOI22_X1 port map( A1 => n6392, A2 => n5064, B1 => n6393, B2 => 
                           n5065, ZN => n6466);
   U6982 : NAND3_X1 port map( A1 => n6470, A2 => n6471, A3 => n6472, ZN => 
                           n12876);
   U6983 : AOI221_X1 port map( B1 => n6385, B2 => n5069, C1 => n6386, C2 => 
                           MEM_IN(20), A => n6473, ZN => n6472);
   U6984 : OAI22_X1 port map( A1 => n11513, A2 => n226, B1 => n5071, B2 => 
                           n6389, ZN => n6473);
   U6985 : AOI22_X1 port map( A1 => n6390, A2 => n5072, B1 => n6391, B2 => 
                           n5073, ZN => n6471);
   U6986 : AOI22_X1 port map( A1 => n6392, A2 => n5074, B1 => n6393, B2 => 
                           n5075, ZN => n6470);
   U6987 : NAND3_X1 port map( A1 => n6474, A2 => n6475, A3 => n6476, ZN => 
                           n12875);
   U6988 : AOI221_X1 port map( B1 => n6385, B2 => n5079, C1 => n6386, C2 => 
                           MEM_IN(21), A => n6477, ZN => n6476);
   U6989 : OAI22_X1 port map( A1 => n11512, A2 => n226, B1 => n5081, B2 => 
                           n6389, ZN => n6477);
   U6990 : AOI22_X1 port map( A1 => n6390, A2 => n5082, B1 => n6391, B2 => 
                           n5083, ZN => n6475);
   U6991 : AOI22_X1 port map( A1 => n6392, A2 => n5084, B1 => n6393, B2 => 
                           n5085, ZN => n6474);
   U6992 : NAND3_X1 port map( A1 => n6478, A2 => n6479, A3 => n6480, ZN => 
                           n12874);
   U6993 : AOI221_X1 port map( B1 => n6385, B2 => n5089, C1 => n6386, C2 => 
                           MEM_IN(22), A => n6481, ZN => n6480);
   U6994 : OAI22_X1 port map( A1 => n11511, A2 => n226, B1 => n5091, B2 => 
                           n6389, ZN => n6481);
   U6995 : AOI22_X1 port map( A1 => n6390, A2 => n5092, B1 => n6391, B2 => 
                           n5093, ZN => n6479);
   U6996 : AOI22_X1 port map( A1 => n6392, A2 => n5094, B1 => n6393, B2 => 
                           n5095, ZN => n6478);
   U6997 : NAND3_X1 port map( A1 => n6482, A2 => n6483, A3 => n6484, ZN => 
                           n12873);
   U6998 : AOI221_X1 port map( B1 => n6385, B2 => n5099, C1 => n6386, C2 => 
                           MEM_IN(23), A => n6485, ZN => n6484);
   U6999 : OAI22_X1 port map( A1 => n11510, A2 => n226, B1 => n5101, B2 => 
                           n6389, ZN => n6485);
   U7000 : AOI22_X1 port map( A1 => n6390, A2 => n5102, B1 => n6391, B2 => 
                           n5103, ZN => n6483);
   U7001 : AOI22_X1 port map( A1 => n6392, A2 => n5104, B1 => n6393, B2 => 
                           n5105, ZN => n6482);
   U7002 : NAND3_X1 port map( A1 => n6486, A2 => n6487, A3 => n6488, ZN => 
                           n12872);
   U7003 : AOI221_X1 port map( B1 => n6385, B2 => n5109, C1 => n6386, C2 => 
                           MEM_IN(24), A => n6489, ZN => n6488);
   U7004 : OAI22_X1 port map( A1 => n11509, A2 => n226, B1 => n5111, B2 => 
                           n6389, ZN => n6489);
   U7005 : AOI22_X1 port map( A1 => n6390, A2 => n5112, B1 => n6391, B2 => 
                           n5113, ZN => n6487);
   U7006 : AOI22_X1 port map( A1 => n6392, A2 => n5114, B1 => n6393, B2 => 
                           n5115, ZN => n6486);
   U7007 : NAND3_X1 port map( A1 => n6490, A2 => n6491, A3 => n6492, ZN => 
                           n12871);
   U7008 : AOI221_X1 port map( B1 => n6385, B2 => n5119, C1 => n6386, C2 => 
                           MEM_IN(25), A => n6493, ZN => n6492);
   U7009 : OAI22_X1 port map( A1 => n11508, A2 => n226, B1 => n5121, B2 => 
                           n6389, ZN => n6493);
   U7010 : AOI22_X1 port map( A1 => n6390, A2 => n5122, B1 => n6391, B2 => 
                           n5123, ZN => n6491);
   U7011 : AOI22_X1 port map( A1 => n6392, A2 => n5124, B1 => n6393, B2 => 
                           n5125, ZN => n6490);
   U7012 : NAND3_X1 port map( A1 => n6494, A2 => n6495, A3 => n6496, ZN => 
                           n12870);
   U7013 : AOI221_X1 port map( B1 => n6385, B2 => n5129, C1 => n6386, C2 => 
                           MEM_IN(26), A => n6497, ZN => n6496);
   U7014 : OAI22_X1 port map( A1 => n11507, A2 => n226, B1 => n5131, B2 => 
                           n6389, ZN => n6497);
   U7015 : AOI22_X1 port map( A1 => n6390, A2 => n5132, B1 => n6391, B2 => 
                           n5133, ZN => n6495);
   U7016 : AOI22_X1 port map( A1 => n6392, A2 => n5134, B1 => n6393, B2 => 
                           n5135, ZN => n6494);
   U7017 : NAND3_X1 port map( A1 => n6498, A2 => n6499, A3 => n6500, ZN => 
                           n12869);
   U7018 : AOI221_X1 port map( B1 => n6385, B2 => n5139, C1 => n6386, C2 => 
                           MEM_IN(27), A => n6501, ZN => n6500);
   U7019 : OAI22_X1 port map( A1 => n11506, A2 => n226, B1 => n5141, B2 => 
                           n6389, ZN => n6501);
   U7020 : AOI22_X1 port map( A1 => n6390, A2 => n5142, B1 => n6391, B2 => 
                           n5143, ZN => n6499);
   U7021 : AOI22_X1 port map( A1 => n6392, A2 => n5144, B1 => n6393, B2 => 
                           n5145, ZN => n6498);
   U7022 : NAND3_X1 port map( A1 => n6502, A2 => n6503, A3 => n6504, ZN => 
                           n12868);
   U7023 : AOI221_X1 port map( B1 => n6385, B2 => n5149, C1 => n6386, C2 => 
                           MEM_IN(28), A => n6505, ZN => n6504);
   U7024 : OAI22_X1 port map( A1 => n11505, A2 => n226, B1 => n5151, B2 => 
                           n6389, ZN => n6505);
   U7025 : AOI22_X1 port map( A1 => n6390, A2 => n5152, B1 => n6391, B2 => 
                           n5153, ZN => n6503);
   U7026 : AOI22_X1 port map( A1 => n6392, A2 => n5154, B1 => n6393, B2 => 
                           n5155, ZN => n6502);
   U7027 : NAND3_X1 port map( A1 => n6506, A2 => n6507, A3 => n6508, ZN => 
                           n12867);
   U7028 : AOI221_X1 port map( B1 => n6385, B2 => n5159, C1 => n6386, C2 => 
                           MEM_IN(29), A => n6509, ZN => n6508);
   U7029 : OAI22_X1 port map( A1 => n11504, A2 => n226, B1 => n5161, B2 => 
                           n6389, ZN => n6509);
   U7030 : AOI22_X1 port map( A1 => n6390, A2 => n5162, B1 => n6391, B2 => 
                           n5163, ZN => n6507);
   U7031 : AOI22_X1 port map( A1 => n6392, A2 => n5164, B1 => n6393, B2 => 
                           n5165, ZN => n6506);
   U7032 : NAND3_X1 port map( A1 => n6510, A2 => n6511, A3 => n6512, ZN => 
                           n12866);
   U7033 : AOI221_X1 port map( B1 => n6385, B2 => n5169, C1 => n6386, C2 => 
                           MEM_IN(30), A => n6513, ZN => n6512);
   U7034 : OAI22_X1 port map( A1 => n11503, A2 => n226, B1 => n5171, B2 => 
                           n6389, ZN => n6513);
   U7035 : AOI22_X1 port map( A1 => n6390, A2 => n5172, B1 => n6391, B2 => 
                           n5173, ZN => n6511);
   U7036 : AOI22_X1 port map( A1 => n6392, A2 => n5174, B1 => n6393, B2 => 
                           n5175, ZN => n6510);
   U7037 : NAND3_X1 port map( A1 => n6514, A2 => n6515, A3 => n6516, ZN => 
                           n12865);
   U7038 : AOI221_X1 port map( B1 => n6385, B2 => n5179, C1 => n6386, C2 => 
                           MEM_IN(31), A => n6517, ZN => n6516);
   U7039 : OAI22_X1 port map( A1 => n11502, A2 => n226, B1 => n5181, B2 => 
                           n6389, ZN => n6517);
   U7040 : INV_X1 port map( A => n6069, ZN => n6066);
   U7041 : AOI22_X1 port map( A1 => n6390, A2 => n5191, B1 => n6391, B2 => 
                           n5192, ZN => n6515);
   U7042 : AOI22_X1 port map( A1 => n6392, A2 => n5195, B1 => n6393, B2 => 
                           n5196, ZN => n6514);
   U7043 : OAI22_X1 port map( A1 => n6519, A2 => n6523, B1 => n208, B2 => n225,
                           ZN => n6520);
   U7044 : INV_X1 port map( A => n6518, ZN => n6523);
   U7045 : NOR3_X1 port map( A1 => n4841, A2 => n225, A3 => n5370, ZN => n6518)
                           ;
   U7046 : OAI22_X1 port map( A1 => n4786, A2 => n6524, B1 => n6525, B2 => 
                           n5204, ZN => n6388);
   U7047 : NOR2_X1 port map( A1 => n5370, A2 => n6519, ZN => n6525);
   U7048 : NAND3_X1 port map( A1 => n6222, A2 => n6225, A3 => n6526, ZN => 
                           n5370);
   U7049 : AOI211_X1 port map( C1 => n6527, C2 => n5207, A => n6528, B => n6069
                           , ZN => n6524);
   U7050 : NAND2_X1 port map( A1 => n6529, A2 => n6530, ZN => n6519);
   U7051 : NOR2_X1 port map( A1 => n6225, A2 => n4787, ZN => n6069);
   U7052 : NAND2_X1 port map( A1 => n6531, A2 => n5215, ZN => n6225);
   U7053 : NAND3_X1 port map( A1 => n6532, A2 => n6533, A3 => n6534, ZN => 
                           n12864);
   U7054 : AOI221_X1 port map( B1 => n6535, B2 => n4863, C1 => n6536, C2 => 
                           MEM_IN(0), A => n6537, ZN => n6534);
   U7055 : OAI22_X1 port map( A1 => n11501, A2 => n228, B1 => n4867, B2 => 
                           n6539, ZN => n6537);
   U7056 : AOI22_X1 port map( A1 => n6540, A2 => n4869, B1 => n6541, B2 => 
                           n4871, ZN => n6533);
   U7057 : AOI22_X1 port map( A1 => n6542, A2 => n4873, B1 => n6543, B2 => 
                           n4875, ZN => n6532);
   U7058 : NAND3_X1 port map( A1 => n6544, A2 => n6545, A3 => n6546, ZN => 
                           n12863);
   U7059 : AOI221_X1 port map( B1 => n6535, B2 => n4879, C1 => n6536, C2 => 
                           MEM_IN(1), A => n6547, ZN => n6546);
   U7060 : OAI22_X1 port map( A1 => n11500, A2 => n228, B1 => n4881, B2 => 
                           n6539, ZN => n6547);
   U7061 : AOI22_X1 port map( A1 => n6540, A2 => n4882, B1 => n6541, B2 => 
                           n4883, ZN => n6545);
   U7062 : AOI22_X1 port map( A1 => n6542, A2 => n4884, B1 => n6543, B2 => 
                           n4885, ZN => n6544);
   U7063 : NAND3_X1 port map( A1 => n6548, A2 => n6549, A3 => n6550, ZN => 
                           n12862);
   U7064 : AOI221_X1 port map( B1 => n6535, B2 => n4889, C1 => n6536, C2 => 
                           MEM_IN(2), A => n6551, ZN => n6550);
   U7065 : OAI22_X1 port map( A1 => n11499, A2 => n228, B1 => n4891, B2 => 
                           n6539, ZN => n6551);
   U7066 : AOI22_X1 port map( A1 => n6540, A2 => n4892, B1 => n6541, B2 => 
                           n4893, ZN => n6549);
   U7067 : AOI22_X1 port map( A1 => n6542, A2 => n4894, B1 => n6543, B2 => 
                           n4895, ZN => n6548);
   U7068 : NAND3_X1 port map( A1 => n6552, A2 => n6553, A3 => n6554, ZN => 
                           n12861);
   U7069 : AOI221_X1 port map( B1 => n6535, B2 => n4899, C1 => n6536, C2 => 
                           MEM_IN(3), A => n6555, ZN => n6554);
   U7070 : OAI22_X1 port map( A1 => n11498, A2 => n228, B1 => n4901, B2 => 
                           n6539, ZN => n6555);
   U7071 : AOI22_X1 port map( A1 => n6540, A2 => n4902, B1 => n6541, B2 => 
                           n4903, ZN => n6553);
   U7072 : AOI22_X1 port map( A1 => n6542, A2 => n4904, B1 => n6543, B2 => 
                           n4905, ZN => n6552);
   U7073 : NAND3_X1 port map( A1 => n6556, A2 => n6557, A3 => n6558, ZN => 
                           n12860);
   U7074 : AOI221_X1 port map( B1 => n6535, B2 => n4909, C1 => n6536, C2 => 
                           MEM_IN(4), A => n6559, ZN => n6558);
   U7075 : OAI22_X1 port map( A1 => n11497, A2 => n228, B1 => n4911, B2 => 
                           n6539, ZN => n6559);
   U7076 : AOI22_X1 port map( A1 => n6540, A2 => n4912, B1 => n6541, B2 => 
                           n4913, ZN => n6557);
   U7077 : AOI22_X1 port map( A1 => n6542, A2 => n4914, B1 => n6543, B2 => 
                           n4915, ZN => n6556);
   U7078 : NAND3_X1 port map( A1 => n6560, A2 => n6561, A3 => n6562, ZN => 
                           n12859);
   U7079 : AOI221_X1 port map( B1 => n6535, B2 => n4919, C1 => n6536, C2 => 
                           MEM_IN(5), A => n6563, ZN => n6562);
   U7080 : OAI22_X1 port map( A1 => n11496, A2 => n228, B1 => n4921, B2 => 
                           n6539, ZN => n6563);
   U7081 : AOI22_X1 port map( A1 => n6540, A2 => n4922, B1 => n6541, B2 => 
                           n4923, ZN => n6561);
   U7082 : AOI22_X1 port map( A1 => n6542, A2 => n4924, B1 => n6543, B2 => 
                           n4925, ZN => n6560);
   U7083 : NAND3_X1 port map( A1 => n6564, A2 => n6565, A3 => n6566, ZN => 
                           n12858);
   U7084 : AOI221_X1 port map( B1 => n6535, B2 => n4929, C1 => n6536, C2 => 
                           MEM_IN(6), A => n6567, ZN => n6566);
   U7085 : OAI22_X1 port map( A1 => n11495, A2 => n228, B1 => n4931, B2 => 
                           n6539, ZN => n6567);
   U7086 : AOI22_X1 port map( A1 => n6540, A2 => n4932, B1 => n6541, B2 => 
                           n4933, ZN => n6565);
   U7087 : AOI22_X1 port map( A1 => n6542, A2 => n4934, B1 => n6543, B2 => 
                           n4935, ZN => n6564);
   U7088 : NAND3_X1 port map( A1 => n6568, A2 => n6569, A3 => n6570, ZN => 
                           n12857);
   U7089 : AOI221_X1 port map( B1 => n6535, B2 => n4939, C1 => n6536, C2 => 
                           MEM_IN(7), A => n6571, ZN => n6570);
   U7090 : OAI22_X1 port map( A1 => n11494, A2 => n228, B1 => n4941, B2 => 
                           n6539, ZN => n6571);
   U7091 : AOI22_X1 port map( A1 => n6540, A2 => n4942, B1 => n6541, B2 => 
                           n4943, ZN => n6569);
   U7092 : AOI22_X1 port map( A1 => n6542, A2 => n4944, B1 => n6543, B2 => 
                           n4945, ZN => n6568);
   U7093 : NAND3_X1 port map( A1 => n6572, A2 => n6573, A3 => n6574, ZN => 
                           n12856);
   U7094 : AOI221_X1 port map( B1 => n6535, B2 => n4949, C1 => n6536, C2 => 
                           MEM_IN(8), A => n6575, ZN => n6574);
   U7095 : OAI22_X1 port map( A1 => n11493, A2 => n228, B1 => n4951, B2 => 
                           n6539, ZN => n6575);
   U7096 : AOI22_X1 port map( A1 => n6540, A2 => n4952, B1 => n6541, B2 => 
                           n4953, ZN => n6573);
   U7097 : AOI22_X1 port map( A1 => n6542, A2 => n4954, B1 => n6543, B2 => 
                           n4955, ZN => n6572);
   U7098 : NAND3_X1 port map( A1 => n6576, A2 => n6577, A3 => n6578, ZN => 
                           n12855);
   U7099 : AOI221_X1 port map( B1 => n6535, B2 => n4959, C1 => n6536, C2 => 
                           MEM_IN(9), A => n6579, ZN => n6578);
   U7100 : OAI22_X1 port map( A1 => n11492, A2 => n228, B1 => n4961, B2 => 
                           n6539, ZN => n6579);
   U7101 : AOI22_X1 port map( A1 => n6540, A2 => n4962, B1 => n6541, B2 => 
                           n4963, ZN => n6577);
   U7102 : AOI22_X1 port map( A1 => n6542, A2 => n4964, B1 => n6543, B2 => 
                           n4965, ZN => n6576);
   U7103 : NAND3_X1 port map( A1 => n6580, A2 => n6581, A3 => n6582, ZN => 
                           n12854);
   U7104 : AOI221_X1 port map( B1 => n6535, B2 => n4969, C1 => n6536, C2 => 
                           MEM_IN(10), A => n6583, ZN => n6582);
   U7105 : OAI22_X1 port map( A1 => n11491, A2 => n228, B1 => n4971, B2 => 
                           n6539, ZN => n6583);
   U7106 : AOI22_X1 port map( A1 => n6540, A2 => n4972, B1 => n6541, B2 => 
                           n4973, ZN => n6581);
   U7107 : AOI22_X1 port map( A1 => n6542, A2 => n4974, B1 => n6543, B2 => 
                           n4975, ZN => n6580);
   U7108 : NAND3_X1 port map( A1 => n6584, A2 => n6585, A3 => n6586, ZN => 
                           n12853);
   U7109 : AOI221_X1 port map( B1 => n6535, B2 => n4979, C1 => n6536, C2 => 
                           MEM_IN(11), A => n6587, ZN => n6586);
   U7110 : OAI22_X1 port map( A1 => n11490, A2 => n228, B1 => n4981, B2 => 
                           n6539, ZN => n6587);
   U7111 : AOI22_X1 port map( A1 => n6540, A2 => n4982, B1 => n6541, B2 => 
                           n4983, ZN => n6585);
   U7112 : AOI22_X1 port map( A1 => n6542, A2 => n4984, B1 => n6543, B2 => 
                           n4985, ZN => n6584);
   U7113 : NAND3_X1 port map( A1 => n6588, A2 => n6589, A3 => n6590, ZN => 
                           n12852);
   U7114 : AOI221_X1 port map( B1 => n6535, B2 => n4989, C1 => n6536, C2 => 
                           MEM_IN(12), A => n6591, ZN => n6590);
   U7115 : OAI22_X1 port map( A1 => n11489, A2 => n228, B1 => n4991, B2 => 
                           n6539, ZN => n6591);
   U7116 : AOI22_X1 port map( A1 => n6540, A2 => n4992, B1 => n6541, B2 => 
                           n4993, ZN => n6589);
   U7117 : AOI22_X1 port map( A1 => n6542, A2 => n4994, B1 => n6543, B2 => 
                           n4995, ZN => n6588);
   U7118 : NAND3_X1 port map( A1 => n6592, A2 => n6593, A3 => n6594, ZN => 
                           n12851);
   U7119 : AOI221_X1 port map( B1 => n6535, B2 => n4999, C1 => n6536, C2 => 
                           MEM_IN(13), A => n6595, ZN => n6594);
   U7120 : OAI22_X1 port map( A1 => n11488, A2 => n228, B1 => n5001, B2 => 
                           n6539, ZN => n6595);
   U7121 : AOI22_X1 port map( A1 => n6540, A2 => n5002, B1 => n6541, B2 => 
                           n5003, ZN => n6593);
   U7122 : AOI22_X1 port map( A1 => n6542, A2 => n5004, B1 => n6543, B2 => 
                           n5005, ZN => n6592);
   U7123 : NAND3_X1 port map( A1 => n6596, A2 => n6597, A3 => n6598, ZN => 
                           n12850);
   U7124 : AOI221_X1 port map( B1 => n6535, B2 => n5009, C1 => n6536, C2 => 
                           MEM_IN(14), A => n6599, ZN => n6598);
   U7125 : OAI22_X1 port map( A1 => n11487, A2 => n228, B1 => n5011, B2 => 
                           n6539, ZN => n6599);
   U7126 : AOI22_X1 port map( A1 => n6540, A2 => n5012, B1 => n6541, B2 => 
                           n5013, ZN => n6597);
   U7127 : AOI22_X1 port map( A1 => n6542, A2 => n5014, B1 => n6543, B2 => 
                           n5015, ZN => n6596);
   U7128 : NAND3_X1 port map( A1 => n6600, A2 => n6601, A3 => n6602, ZN => 
                           n12849);
   U7129 : AOI221_X1 port map( B1 => n6535, B2 => n5019, C1 => n6536, C2 => 
                           MEM_IN(15), A => n6603, ZN => n6602);
   U7130 : OAI22_X1 port map( A1 => n11486, A2 => n228, B1 => n5021, B2 => 
                           n6539, ZN => n6603);
   U7131 : AOI22_X1 port map( A1 => n6540, A2 => n5022, B1 => n6541, B2 => 
                           n5023, ZN => n6601);
   U7132 : AOI22_X1 port map( A1 => n6542, A2 => n5024, B1 => n6543, B2 => 
                           n5025, ZN => n6600);
   U7133 : NAND3_X1 port map( A1 => n6604, A2 => n6605, A3 => n6606, ZN => 
                           n12848);
   U7134 : AOI221_X1 port map( B1 => n6535, B2 => n5029, C1 => n6536, C2 => 
                           MEM_IN(16), A => n6607, ZN => n6606);
   U7135 : OAI22_X1 port map( A1 => n11485, A2 => n228, B1 => n5031, B2 => 
                           n6539, ZN => n6607);
   U7136 : AOI22_X1 port map( A1 => n6540, A2 => n5032, B1 => n6541, B2 => 
                           n5033, ZN => n6605);
   U7137 : AOI22_X1 port map( A1 => n6542, A2 => n5034, B1 => n6543, B2 => 
                           n5035, ZN => n6604);
   U7138 : NAND3_X1 port map( A1 => n6608, A2 => n6609, A3 => n6610, ZN => 
                           n12847);
   U7139 : AOI221_X1 port map( B1 => n6535, B2 => n5039, C1 => n6536, C2 => 
                           MEM_IN(17), A => n6611, ZN => n6610);
   U7140 : OAI22_X1 port map( A1 => n11484, A2 => n228, B1 => n5041, B2 => 
                           n6539, ZN => n6611);
   U7141 : AOI22_X1 port map( A1 => n6540, A2 => n5042, B1 => n6541, B2 => 
                           n5043, ZN => n6609);
   U7142 : AOI22_X1 port map( A1 => n6542, A2 => n5044, B1 => n6543, B2 => 
                           n5045, ZN => n6608);
   U7143 : NAND3_X1 port map( A1 => n6612, A2 => n6613, A3 => n6614, ZN => 
                           n12846);
   U7144 : AOI221_X1 port map( B1 => n6535, B2 => n5049, C1 => n6536, C2 => 
                           MEM_IN(18), A => n6615, ZN => n6614);
   U7145 : OAI22_X1 port map( A1 => n11483, A2 => n228, B1 => n5051, B2 => 
                           n6539, ZN => n6615);
   U7146 : AOI22_X1 port map( A1 => n6540, A2 => n5052, B1 => n6541, B2 => 
                           n5053, ZN => n6613);
   U7147 : AOI22_X1 port map( A1 => n6542, A2 => n5054, B1 => n6543, B2 => 
                           n5055, ZN => n6612);
   U7148 : NAND3_X1 port map( A1 => n6616, A2 => n6617, A3 => n6618, ZN => 
                           n12845);
   U7149 : AOI221_X1 port map( B1 => n6535, B2 => n5059, C1 => n6536, C2 => 
                           MEM_IN(19), A => n6619, ZN => n6618);
   U7150 : OAI22_X1 port map( A1 => n11482, A2 => n228, B1 => n5061, B2 => 
                           n6539, ZN => n6619);
   U7151 : AOI22_X1 port map( A1 => n6540, A2 => n5062, B1 => n6541, B2 => 
                           n5063, ZN => n6617);
   U7152 : AOI22_X1 port map( A1 => n6542, A2 => n5064, B1 => n6543, B2 => 
                           n5065, ZN => n6616);
   U7153 : NAND3_X1 port map( A1 => n6620, A2 => n6621, A3 => n6622, ZN => 
                           n12844);
   U7154 : AOI221_X1 port map( B1 => n6535, B2 => n5069, C1 => n6536, C2 => 
                           MEM_IN(20), A => n6623, ZN => n6622);
   U7155 : OAI22_X1 port map( A1 => n11481, A2 => n228, B1 => n5071, B2 => 
                           n6539, ZN => n6623);
   U7156 : AOI22_X1 port map( A1 => n6540, A2 => n5072, B1 => n6541, B2 => 
                           n5073, ZN => n6621);
   U7157 : AOI22_X1 port map( A1 => n6542, A2 => n5074, B1 => n6543, B2 => 
                           n5075, ZN => n6620);
   U7158 : NAND3_X1 port map( A1 => n6624, A2 => n6625, A3 => n6626, ZN => 
                           n12843);
   U7159 : AOI221_X1 port map( B1 => n6535, B2 => n5079, C1 => n6536, C2 => 
                           MEM_IN(21), A => n6627, ZN => n6626);
   U7160 : OAI22_X1 port map( A1 => n11480, A2 => n228, B1 => n5081, B2 => 
                           n6539, ZN => n6627);
   U7161 : AOI22_X1 port map( A1 => n6540, A2 => n5082, B1 => n6541, B2 => 
                           n5083, ZN => n6625);
   U7162 : AOI22_X1 port map( A1 => n6542, A2 => n5084, B1 => n6543, B2 => 
                           n5085, ZN => n6624);
   U7163 : NAND3_X1 port map( A1 => n6628, A2 => n6629, A3 => n6630, ZN => 
                           n12842);
   U7164 : AOI221_X1 port map( B1 => n6535, B2 => n5089, C1 => n6536, C2 => 
                           MEM_IN(22), A => n6631, ZN => n6630);
   U7165 : OAI22_X1 port map( A1 => n11479, A2 => n228, B1 => n5091, B2 => 
                           n6539, ZN => n6631);
   U7166 : AOI22_X1 port map( A1 => n6540, A2 => n5092, B1 => n6541, B2 => 
                           n5093, ZN => n6629);
   U7167 : AOI22_X1 port map( A1 => n6542, A2 => n5094, B1 => n6543, B2 => 
                           n5095, ZN => n6628);
   U7168 : NAND3_X1 port map( A1 => n6632, A2 => n6633, A3 => n6634, ZN => 
                           n12841);
   U7169 : AOI221_X1 port map( B1 => n6535, B2 => n5099, C1 => n6536, C2 => 
                           MEM_IN(23), A => n6635, ZN => n6634);
   U7170 : OAI22_X1 port map( A1 => n11478, A2 => n228, B1 => n5101, B2 => 
                           n6539, ZN => n6635);
   U7171 : AOI22_X1 port map( A1 => n6540, A2 => n5102, B1 => n6541, B2 => 
                           n5103, ZN => n6633);
   U7172 : AOI22_X1 port map( A1 => n6542, A2 => n5104, B1 => n6543, B2 => 
                           n5105, ZN => n6632);
   U7173 : NAND3_X1 port map( A1 => n6636, A2 => n6637, A3 => n6638, ZN => 
                           n12840);
   U7174 : AOI221_X1 port map( B1 => n6535, B2 => n5109, C1 => n6536, C2 => 
                           MEM_IN(24), A => n6639, ZN => n6638);
   U7175 : OAI22_X1 port map( A1 => n11477, A2 => n228, B1 => n5111, B2 => 
                           n6539, ZN => n6639);
   U7176 : AOI22_X1 port map( A1 => n6540, A2 => n5112, B1 => n6541, B2 => 
                           n5113, ZN => n6637);
   U7177 : AOI22_X1 port map( A1 => n6542, A2 => n5114, B1 => n6543, B2 => 
                           n5115, ZN => n6636);
   U7178 : NAND3_X1 port map( A1 => n6640, A2 => n6641, A3 => n6642, ZN => 
                           n12839);
   U7179 : AOI221_X1 port map( B1 => n6535, B2 => n5119, C1 => n6536, C2 => 
                           MEM_IN(25), A => n6643, ZN => n6642);
   U7180 : OAI22_X1 port map( A1 => n11476, A2 => n228, B1 => n5121, B2 => 
                           n6539, ZN => n6643);
   U7181 : AOI22_X1 port map( A1 => n6540, A2 => n5122, B1 => n6541, B2 => 
                           n5123, ZN => n6641);
   U7182 : AOI22_X1 port map( A1 => n6542, A2 => n5124, B1 => n6543, B2 => 
                           n5125, ZN => n6640);
   U7183 : NAND3_X1 port map( A1 => n6644, A2 => n6645, A3 => n6646, ZN => 
                           n12838);
   U7184 : AOI221_X1 port map( B1 => n6535, B2 => n5129, C1 => n6536, C2 => 
                           MEM_IN(26), A => n6647, ZN => n6646);
   U7185 : OAI22_X1 port map( A1 => n11475, A2 => n228, B1 => n5131, B2 => 
                           n6539, ZN => n6647);
   U7186 : AOI22_X1 port map( A1 => n6540, A2 => n5132, B1 => n6541, B2 => 
                           n5133, ZN => n6645);
   U7187 : AOI22_X1 port map( A1 => n6542, A2 => n5134, B1 => n6543, B2 => 
                           n5135, ZN => n6644);
   U7188 : NAND3_X1 port map( A1 => n6648, A2 => n6649, A3 => n6650, ZN => 
                           n12837);
   U7189 : AOI221_X1 port map( B1 => n6535, B2 => n5139, C1 => n6536, C2 => 
                           MEM_IN(27), A => n6651, ZN => n6650);
   U7190 : OAI22_X1 port map( A1 => n11474, A2 => n228, B1 => n5141, B2 => 
                           n6539, ZN => n6651);
   U7191 : AOI22_X1 port map( A1 => n6540, A2 => n5142, B1 => n6541, B2 => 
                           n5143, ZN => n6649);
   U7192 : AOI22_X1 port map( A1 => n6542, A2 => n5144, B1 => n6543, B2 => 
                           n5145, ZN => n6648);
   U7193 : NAND3_X1 port map( A1 => n6652, A2 => n6653, A3 => n6654, ZN => 
                           n12836);
   U7194 : AOI221_X1 port map( B1 => n6535, B2 => n5149, C1 => n6536, C2 => 
                           MEM_IN(28), A => n6655, ZN => n6654);
   U7195 : OAI22_X1 port map( A1 => n11473, A2 => n228, B1 => n5151, B2 => 
                           n6539, ZN => n6655);
   U7196 : AOI22_X1 port map( A1 => n6540, A2 => n5152, B1 => n6541, B2 => 
                           n5153, ZN => n6653);
   U7197 : AOI22_X1 port map( A1 => n6542, A2 => n5154, B1 => n6543, B2 => 
                           n5155, ZN => n6652);
   U7198 : NAND3_X1 port map( A1 => n6656, A2 => n6657, A3 => n6658, ZN => 
                           n12835);
   U7199 : AOI221_X1 port map( B1 => n6535, B2 => n5159, C1 => n6536, C2 => 
                           MEM_IN(29), A => n6659, ZN => n6658);
   U7200 : OAI22_X1 port map( A1 => n11472, A2 => n228, B1 => n5161, B2 => 
                           n6539, ZN => n6659);
   U7201 : AOI22_X1 port map( A1 => n6540, A2 => n5162, B1 => n6541, B2 => 
                           n5163, ZN => n6657);
   U7202 : AOI22_X1 port map( A1 => n6542, A2 => n5164, B1 => n6543, B2 => 
                           n5165, ZN => n6656);
   U7203 : NAND3_X1 port map( A1 => n6660, A2 => n6661, A3 => n6662, ZN => 
                           n12834);
   U7204 : AOI221_X1 port map( B1 => n6535, B2 => n5169, C1 => n6536, C2 => 
                           MEM_IN(30), A => n6663, ZN => n6662);
   U7205 : OAI22_X1 port map( A1 => n11471, A2 => n228, B1 => n5171, B2 => 
                           n6539, ZN => n6663);
   U7206 : AOI22_X1 port map( A1 => n6540, A2 => n5172, B1 => n6541, B2 => 
                           n5173, ZN => n6661);
   U7207 : AOI22_X1 port map( A1 => n6542, A2 => n5174, B1 => n6543, B2 => 
                           n5175, ZN => n6660);
   U7208 : NAND3_X1 port map( A1 => n6664, A2 => n6665, A3 => n6666, ZN => 
                           n12833);
   U7209 : AOI221_X1 port map( B1 => n6535, B2 => n5179, C1 => n6536, C2 => 
                           MEM_IN(31), A => n6667, ZN => n6666);
   U7210 : OAI22_X1 port map( A1 => n11470, A2 => n228, B1 => n5181, B2 => 
                           n6539, ZN => n6667);
   U7211 : NAND2_X1 port map( A1 => n5206, A2 => n6074, ZN => n6368);
   U7212 : AOI22_X1 port map( A1 => n6540, A2 => n5191, B1 => n6541, B2 => 
                           n5192, ZN => n6665);
   U7213 : AOI22_X1 port map( A1 => n6542, A2 => n5195, B1 => n6543, B2 => 
                           n5196, ZN => n6664);
   U7214 : OAI22_X1 port map( A1 => n6669, A2 => n6673, B1 => n208, B2 => n227,
                           ZN => n6670);
   U7215 : INV_X1 port map( A => n6668, ZN => n6673);
   U7216 : NOR3_X1 port map( A1 => n4841, A2 => n227, A3 => n5524, ZN => n6668)
                           ;
   U7217 : OAI22_X1 port map( A1 => n4786, A2 => n6674, B1 => n6675, B2 => 
                           n5204, ZN => n6538);
   U7218 : NOR2_X1 port map( A1 => n5524, A2 => n6669, ZN => n6675);
   U7219 : NAND2_X1 port map( A1 => n6676, A2 => n6222, ZN => n5524);
   U7220 : AOI211_X1 port map( C1 => n6527, C2 => n5365, A => n6528, B => n6672
                           , ZN => n6674);
   U7221 : OAI21_X1 port map( B1 => n6222, B2 => n4787, A => n5368, ZN => n6528
                           );
   U7222 : NOR2_X1 port map( A1 => n6074, A2 => n6078, ZN => n6222);
   U7223 : NAND2_X1 port map( A1 => n5925, A2 => n5774, ZN => n6074);
   U7224 : NAND2_X1 port map( A1 => n6677, A2 => n6678, ZN => n6669);
   U7225 : NOR2_X1 port map( A1 => n5774, A2 => n4787, ZN => n6224);
   U7226 : NAND2_X1 port map( A1 => n6531, A2 => n5372, ZN => n5774);
   U7227 : NAND3_X1 port map( A1 => n6679, A2 => n6680, A3 => n6681, ZN => 
                           n12832);
   U7228 : AOI221_X1 port map( B1 => n219, B2 => n4863, C1 => n6682, C2 => 
                           MEM_IN(0), A => n6683, ZN => n6681);
   U7229 : OAI22_X1 port map( A1 => n11469, A2 => n247, B1 => n4867, B2 => n148
                           , ZN => n6683);
   U7230 : AOI22_X1 port map( A1 => n198, A2 => n4869, B1 => n163, B2 => n4871,
                           ZN => n6680);
   U7231 : AOI22_X1 port map( A1 => n240, A2 => n4873, B1 => n160, B2 => n4875,
                           ZN => n6679);
   U7232 : NAND3_X1 port map( A1 => n6685, A2 => n6686, A3 => n6687, ZN => 
                           n12831);
   U7233 : AOI221_X1 port map( B1 => n219, B2 => n4879, C1 => n6682, C2 => 
                           MEM_IN(1), A => n6688, ZN => n6687);
   U7234 : OAI22_X1 port map( A1 => n11468, A2 => n247, B1 => n4881, B2 => n148
                           , ZN => n6688);
   U7235 : AOI22_X1 port map( A1 => n198, A2 => n4882, B1 => n163, B2 => n4883,
                           ZN => n6686);
   U7236 : AOI22_X1 port map( A1 => n240, A2 => n4884, B1 => n160, B2 => n4885,
                           ZN => n6685);
   U7237 : NAND3_X1 port map( A1 => n6689, A2 => n6690, A3 => n6691, ZN => 
                           n12830);
   U7238 : AOI221_X1 port map( B1 => n219, B2 => n4889, C1 => n6682, C2 => 
                           MEM_IN(2), A => n6692, ZN => n6691);
   U7239 : OAI22_X1 port map( A1 => n11467, A2 => n247, B1 => n4891, B2 => n148
                           , ZN => n6692);
   U7240 : AOI22_X1 port map( A1 => n198, A2 => n4892, B1 => n163, B2 => n4893,
                           ZN => n6690);
   U7241 : AOI22_X1 port map( A1 => n240, A2 => n4894, B1 => n160, B2 => n4895,
                           ZN => n6689);
   U7242 : NAND3_X1 port map( A1 => n6693, A2 => n6694, A3 => n6695, ZN => 
                           n12829);
   U7243 : AOI221_X1 port map( B1 => n219, B2 => n4899, C1 => n6682, C2 => 
                           MEM_IN(3), A => n6696, ZN => n6695);
   U7244 : OAI22_X1 port map( A1 => n11466, A2 => n247, B1 => n4901, B2 => n148
                           , ZN => n6696);
   U7245 : AOI22_X1 port map( A1 => n198, A2 => n4902, B1 => n163, B2 => n4903,
                           ZN => n6694);
   U7246 : AOI22_X1 port map( A1 => n240, A2 => n4904, B1 => n160, B2 => n4905,
                           ZN => n6693);
   U7247 : NAND3_X1 port map( A1 => n6697, A2 => n6698, A3 => n6699, ZN => 
                           n12828);
   U7248 : AOI221_X1 port map( B1 => n219, B2 => n4909, C1 => n6682, C2 => 
                           MEM_IN(4), A => n6700, ZN => n6699);
   U7249 : OAI22_X1 port map( A1 => n11465, A2 => n247, B1 => n4911, B2 => n148
                           , ZN => n6700);
   U7250 : AOI22_X1 port map( A1 => n198, A2 => n4912, B1 => n163, B2 => n4913,
                           ZN => n6698);
   U7251 : AOI22_X1 port map( A1 => n240, A2 => n4914, B1 => n160, B2 => n4915,
                           ZN => n6697);
   U7252 : NAND3_X1 port map( A1 => n6701, A2 => n6702, A3 => n6703, ZN => 
                           n12827);
   U7253 : AOI221_X1 port map( B1 => n219, B2 => n4919, C1 => n6682, C2 => 
                           MEM_IN(5), A => n6704, ZN => n6703);
   U7254 : OAI22_X1 port map( A1 => n11464, A2 => n247, B1 => n4921, B2 => n148
                           , ZN => n6704);
   U7255 : AOI22_X1 port map( A1 => n198, A2 => n4922, B1 => n163, B2 => n4923,
                           ZN => n6702);
   U7256 : AOI22_X1 port map( A1 => n240, A2 => n4924, B1 => n160, B2 => n4925,
                           ZN => n6701);
   U7257 : NAND3_X1 port map( A1 => n6705, A2 => n6706, A3 => n6707, ZN => 
                           n12826);
   U7258 : AOI221_X1 port map( B1 => n219, B2 => n4929, C1 => n6682, C2 => 
                           MEM_IN(6), A => n6708, ZN => n6707);
   U7259 : OAI22_X1 port map( A1 => n11463, A2 => n247, B1 => n4931, B2 => n148
                           , ZN => n6708);
   U7260 : AOI22_X1 port map( A1 => n198, A2 => n4932, B1 => n163, B2 => n4933,
                           ZN => n6706);
   U7261 : AOI22_X1 port map( A1 => n240, A2 => n4934, B1 => n160, B2 => n4935,
                           ZN => n6705);
   U7262 : NAND3_X1 port map( A1 => n6709, A2 => n6710, A3 => n6711, ZN => 
                           n12825);
   U7263 : AOI221_X1 port map( B1 => n219, B2 => n4939, C1 => n6682, C2 => 
                           MEM_IN(7), A => n6712, ZN => n6711);
   U7264 : OAI22_X1 port map( A1 => n11462, A2 => n247, B1 => n4941, B2 => n148
                           , ZN => n6712);
   U7265 : AOI22_X1 port map( A1 => n198, A2 => n4942, B1 => n163, B2 => n4943,
                           ZN => n6710);
   U7266 : AOI22_X1 port map( A1 => n240, A2 => n4944, B1 => n160, B2 => n4945,
                           ZN => n6709);
   U7267 : NAND3_X1 port map( A1 => n6713, A2 => n6714, A3 => n6715, ZN => 
                           n12824);
   U7268 : AOI221_X1 port map( B1 => n219, B2 => n4949, C1 => n6682, C2 => 
                           MEM_IN(8), A => n6716, ZN => n6715);
   U7269 : OAI22_X1 port map( A1 => n11461, A2 => n247, B1 => n4951, B2 => n148
                           , ZN => n6716);
   U7270 : AOI22_X1 port map( A1 => n198, A2 => n4952, B1 => n163, B2 => n4953,
                           ZN => n6714);
   U7271 : AOI22_X1 port map( A1 => n240, A2 => n4954, B1 => n160, B2 => n4955,
                           ZN => n6713);
   U7272 : NAND3_X1 port map( A1 => n6717, A2 => n6718, A3 => n6719, ZN => 
                           n12823);
   U7273 : AOI221_X1 port map( B1 => n219, B2 => n4959, C1 => n6682, C2 => 
                           MEM_IN(9), A => n6720, ZN => n6719);
   U7274 : OAI22_X1 port map( A1 => n11460, A2 => n247, B1 => n4961, B2 => n148
                           , ZN => n6720);
   U7275 : AOI22_X1 port map( A1 => n198, A2 => n4962, B1 => n163, B2 => n4963,
                           ZN => n6718);
   U7276 : AOI22_X1 port map( A1 => n240, A2 => n4964, B1 => n160, B2 => n4965,
                           ZN => n6717);
   U7277 : NAND3_X1 port map( A1 => n6721, A2 => n6722, A3 => n6723, ZN => 
                           n12822);
   U7278 : AOI221_X1 port map( B1 => n219, B2 => n4969, C1 => n6682, C2 => 
                           MEM_IN(10), A => n6724, ZN => n6723);
   U7279 : OAI22_X1 port map( A1 => n11459, A2 => n247, B1 => n4971, B2 => n148
                           , ZN => n6724);
   U7280 : AOI22_X1 port map( A1 => n198, A2 => n4972, B1 => n163, B2 => n4973,
                           ZN => n6722);
   U7281 : AOI22_X1 port map( A1 => n240, A2 => n4974, B1 => n160, B2 => n4975,
                           ZN => n6721);
   U7282 : NAND3_X1 port map( A1 => n6725, A2 => n6726, A3 => n6727, ZN => 
                           n12821);
   U7283 : AOI221_X1 port map( B1 => n219, B2 => n4979, C1 => n6682, C2 => 
                           MEM_IN(11), A => n6728, ZN => n6727);
   U7284 : OAI22_X1 port map( A1 => n11458, A2 => n247, B1 => n4981, B2 => n148
                           , ZN => n6728);
   U7285 : AOI22_X1 port map( A1 => n198, A2 => n4982, B1 => n163, B2 => n4983,
                           ZN => n6726);
   U7286 : AOI22_X1 port map( A1 => n240, A2 => n4984, B1 => n160, B2 => n4985,
                           ZN => n6725);
   U7287 : NAND3_X1 port map( A1 => n6729, A2 => n6730, A3 => n6731, ZN => 
                           n12820);
   U7288 : AOI221_X1 port map( B1 => n219, B2 => n4989, C1 => n6682, C2 => 
                           MEM_IN(12), A => n6732, ZN => n6731);
   U7289 : OAI22_X1 port map( A1 => n11457, A2 => n247, B1 => n4991, B2 => n148
                           , ZN => n6732);
   U7290 : AOI22_X1 port map( A1 => n198, A2 => n4992, B1 => n163, B2 => n4993,
                           ZN => n6730);
   U7291 : AOI22_X1 port map( A1 => n240, A2 => n4994, B1 => n160, B2 => n4995,
                           ZN => n6729);
   U7292 : NAND3_X1 port map( A1 => n6733, A2 => n6734, A3 => n6735, ZN => 
                           n12819);
   U7293 : AOI221_X1 port map( B1 => n219, B2 => n4999, C1 => n6682, C2 => 
                           MEM_IN(13), A => n6736, ZN => n6735);
   U7294 : OAI22_X1 port map( A1 => n11456, A2 => n247, B1 => n5001, B2 => n148
                           , ZN => n6736);
   U7295 : AOI22_X1 port map( A1 => n198, A2 => n5002, B1 => n163, B2 => n5003,
                           ZN => n6734);
   U7296 : AOI22_X1 port map( A1 => n240, A2 => n5004, B1 => n160, B2 => n5005,
                           ZN => n6733);
   U7297 : NAND3_X1 port map( A1 => n6737, A2 => n6738, A3 => n6739, ZN => 
                           n12818);
   U7298 : AOI221_X1 port map( B1 => n219, B2 => n5009, C1 => n6682, C2 => 
                           MEM_IN(14), A => n6740, ZN => n6739);
   U7299 : OAI22_X1 port map( A1 => n11455, A2 => n247, B1 => n5011, B2 => n148
                           , ZN => n6740);
   U7300 : AOI22_X1 port map( A1 => n198, A2 => n5012, B1 => n163, B2 => n5013,
                           ZN => n6738);
   U7301 : AOI22_X1 port map( A1 => n240, A2 => n5014, B1 => n160, B2 => n5015,
                           ZN => n6737);
   U7302 : NAND3_X1 port map( A1 => n6741, A2 => n6742, A3 => n6743, ZN => 
                           n12817);
   U7303 : AOI221_X1 port map( B1 => n219, B2 => n5019, C1 => n6682, C2 => 
                           MEM_IN(15), A => n6744, ZN => n6743);
   U7304 : OAI22_X1 port map( A1 => n11454, A2 => n247, B1 => n5021, B2 => n148
                           , ZN => n6744);
   U7305 : AOI22_X1 port map( A1 => n198, A2 => n5022, B1 => n163, B2 => n5023,
                           ZN => n6742);
   U7306 : AOI22_X1 port map( A1 => n240, A2 => n5024, B1 => n160, B2 => n5025,
                           ZN => n6741);
   U7307 : NAND3_X1 port map( A1 => n6745, A2 => n6746, A3 => n6747, ZN => 
                           n12816);
   U7308 : AOI221_X1 port map( B1 => n219, B2 => n5029, C1 => n6682, C2 => 
                           MEM_IN(16), A => n6748, ZN => n6747);
   U7309 : OAI22_X1 port map( A1 => n11453, A2 => n247, B1 => n5031, B2 => n148
                           , ZN => n6748);
   U7310 : AOI22_X1 port map( A1 => n198, A2 => n5032, B1 => n163, B2 => n5033,
                           ZN => n6746);
   U7311 : AOI22_X1 port map( A1 => n240, A2 => n5034, B1 => n160, B2 => n5035,
                           ZN => n6745);
   U7312 : NAND3_X1 port map( A1 => n6749, A2 => n6750, A3 => n6751, ZN => 
                           n12815);
   U7313 : AOI221_X1 port map( B1 => n219, B2 => n5039, C1 => n6682, C2 => 
                           MEM_IN(17), A => n6752, ZN => n6751);
   U7314 : OAI22_X1 port map( A1 => n11452, A2 => n247, B1 => n5041, B2 => n148
                           , ZN => n6752);
   U7315 : AOI22_X1 port map( A1 => n198, A2 => n5042, B1 => n163, B2 => n5043,
                           ZN => n6750);
   U7316 : AOI22_X1 port map( A1 => n240, A2 => n5044, B1 => n160, B2 => n5045,
                           ZN => n6749);
   U7317 : NAND3_X1 port map( A1 => n6753, A2 => n6754, A3 => n6755, ZN => 
                           n12814);
   U7318 : AOI221_X1 port map( B1 => n219, B2 => n5049, C1 => n6682, C2 => 
                           MEM_IN(18), A => n6756, ZN => n6755);
   U7319 : OAI22_X1 port map( A1 => n11451, A2 => n247, B1 => n5051, B2 => n148
                           , ZN => n6756);
   U7320 : AOI22_X1 port map( A1 => n198, A2 => n5052, B1 => n163, B2 => n5053,
                           ZN => n6754);
   U7321 : AOI22_X1 port map( A1 => n240, A2 => n5054, B1 => n160, B2 => n5055,
                           ZN => n6753);
   U7322 : NAND3_X1 port map( A1 => n6757, A2 => n6758, A3 => n6759, ZN => 
                           n12813);
   U7323 : AOI221_X1 port map( B1 => n219, B2 => n5059, C1 => n6682, C2 => 
                           MEM_IN(19), A => n6760, ZN => n6759);
   U7324 : OAI22_X1 port map( A1 => n11450, A2 => n247, B1 => n5061, B2 => n148
                           , ZN => n6760);
   U7325 : AOI22_X1 port map( A1 => n198, A2 => n5062, B1 => n163, B2 => n5063,
                           ZN => n6758);
   U7326 : AOI22_X1 port map( A1 => n240, A2 => n5064, B1 => n160, B2 => n5065,
                           ZN => n6757);
   U7327 : NAND3_X1 port map( A1 => n6761, A2 => n6762, A3 => n6763, ZN => 
                           n12812);
   U7328 : AOI221_X1 port map( B1 => n219, B2 => n5069, C1 => n6682, C2 => 
                           MEM_IN(20), A => n6764, ZN => n6763);
   U7329 : OAI22_X1 port map( A1 => n11449, A2 => n247, B1 => n5071, B2 => n148
                           , ZN => n6764);
   U7330 : AOI22_X1 port map( A1 => n198, A2 => n5072, B1 => n163, B2 => n5073,
                           ZN => n6762);
   U7331 : AOI22_X1 port map( A1 => n240, A2 => n5074, B1 => n160, B2 => n5075,
                           ZN => n6761);
   U7332 : NAND3_X1 port map( A1 => n6765, A2 => n6766, A3 => n6767, ZN => 
                           n12811);
   U7333 : AOI221_X1 port map( B1 => n219, B2 => n5079, C1 => n6682, C2 => 
                           MEM_IN(21), A => n6768, ZN => n6767);
   U7334 : OAI22_X1 port map( A1 => n11448, A2 => n247, B1 => n5081, B2 => n148
                           , ZN => n6768);
   U7335 : AOI22_X1 port map( A1 => n198, A2 => n5082, B1 => n163, B2 => n5083,
                           ZN => n6766);
   U7336 : AOI22_X1 port map( A1 => n240, A2 => n5084, B1 => n160, B2 => n5085,
                           ZN => n6765);
   U7337 : NAND3_X1 port map( A1 => n6769, A2 => n6770, A3 => n6771, ZN => 
                           n12810);
   U7338 : AOI221_X1 port map( B1 => n219, B2 => n5089, C1 => n6682, C2 => 
                           MEM_IN(22), A => n6772, ZN => n6771);
   U7339 : OAI22_X1 port map( A1 => n11447, A2 => n247, B1 => n5091, B2 => n148
                           , ZN => n6772);
   U7340 : AOI22_X1 port map( A1 => n198, A2 => n5092, B1 => n163, B2 => n5093,
                           ZN => n6770);
   U7341 : AOI22_X1 port map( A1 => n240, A2 => n5094, B1 => n160, B2 => n5095,
                           ZN => n6769);
   U7342 : NAND3_X1 port map( A1 => n6773, A2 => n6774, A3 => n6775, ZN => 
                           n12809);
   U7343 : AOI221_X1 port map( B1 => n219, B2 => n5099, C1 => n6682, C2 => 
                           MEM_IN(23), A => n6776, ZN => n6775);
   U7344 : OAI22_X1 port map( A1 => n11446, A2 => n247, B1 => n5101, B2 => n148
                           , ZN => n6776);
   U7345 : AOI22_X1 port map( A1 => n198, A2 => n5102, B1 => n163, B2 => n5103,
                           ZN => n6774);
   U7346 : AOI22_X1 port map( A1 => n240, A2 => n5104, B1 => n160, B2 => n5105,
                           ZN => n6773);
   U7347 : NAND3_X1 port map( A1 => n6777, A2 => n6778, A3 => n6779, ZN => 
                           n12808);
   U7348 : AOI221_X1 port map( B1 => n219, B2 => n5109, C1 => n6682, C2 => 
                           MEM_IN(24), A => n6780, ZN => n6779);
   U7349 : OAI22_X1 port map( A1 => n11445, A2 => n247, B1 => n5111, B2 => n148
                           , ZN => n6780);
   U7350 : AOI22_X1 port map( A1 => n198, A2 => n5112, B1 => n163, B2 => n5113,
                           ZN => n6778);
   U7351 : AOI22_X1 port map( A1 => n240, A2 => n5114, B1 => n160, B2 => n5115,
                           ZN => n6777);
   U7352 : NAND3_X1 port map( A1 => n6781, A2 => n6782, A3 => n6783, ZN => 
                           n12807);
   U7353 : AOI221_X1 port map( B1 => n219, B2 => n5119, C1 => n6682, C2 => 
                           MEM_IN(25), A => n6784, ZN => n6783);
   U7354 : OAI22_X1 port map( A1 => n11444, A2 => n247, B1 => n5121, B2 => n148
                           , ZN => n6784);
   U7355 : AOI22_X1 port map( A1 => n198, A2 => n5122, B1 => n163, B2 => n5123,
                           ZN => n6782);
   U7356 : AOI22_X1 port map( A1 => n240, A2 => n5124, B1 => n160, B2 => n5125,
                           ZN => n6781);
   U7357 : NAND3_X1 port map( A1 => n6785, A2 => n6786, A3 => n6787, ZN => 
                           n12806);
   U7358 : AOI221_X1 port map( B1 => n219, B2 => n5129, C1 => n6682, C2 => 
                           MEM_IN(26), A => n6788, ZN => n6787);
   U7359 : OAI22_X1 port map( A1 => n11443, A2 => n247, B1 => n5131, B2 => n148
                           , ZN => n6788);
   U7360 : AOI22_X1 port map( A1 => n198, A2 => n5132, B1 => n163, B2 => n5133,
                           ZN => n6786);
   U7361 : AOI22_X1 port map( A1 => n240, A2 => n5134, B1 => n160, B2 => n5135,
                           ZN => n6785);
   U7362 : NAND3_X1 port map( A1 => n6789, A2 => n6790, A3 => n6791, ZN => 
                           n12805);
   U7363 : AOI221_X1 port map( B1 => n219, B2 => n5139, C1 => n6682, C2 => 
                           MEM_IN(27), A => n6792, ZN => n6791);
   U7364 : OAI22_X1 port map( A1 => n11442, A2 => n247, B1 => n5141, B2 => n148
                           , ZN => n6792);
   U7365 : AOI22_X1 port map( A1 => n198, A2 => n5142, B1 => n163, B2 => n5143,
                           ZN => n6790);
   U7366 : AOI22_X1 port map( A1 => n240, A2 => n5144, B1 => n160, B2 => n5145,
                           ZN => n6789);
   U7367 : NAND3_X1 port map( A1 => n6793, A2 => n6794, A3 => n6795, ZN => 
                           n12804);
   U7368 : AOI221_X1 port map( B1 => n219, B2 => n5149, C1 => n6682, C2 => 
                           MEM_IN(28), A => n6796, ZN => n6795);
   U7369 : OAI22_X1 port map( A1 => n11441, A2 => n247, B1 => n5151, B2 => n148
                           , ZN => n6796);
   U7370 : AOI22_X1 port map( A1 => n198, A2 => n5152, B1 => n163, B2 => n5153,
                           ZN => n6794);
   U7371 : AOI22_X1 port map( A1 => n240, A2 => n5154, B1 => n160, B2 => n5155,
                           ZN => n6793);
   U7372 : NAND3_X1 port map( A1 => n6797, A2 => n6798, A3 => n6799, ZN => 
                           n12803);
   U7373 : AOI221_X1 port map( B1 => n219, B2 => n5159, C1 => n6682, C2 => 
                           MEM_IN(29), A => n6800, ZN => n6799);
   U7374 : OAI22_X1 port map( A1 => n11440, A2 => n247, B1 => n5161, B2 => n148
                           , ZN => n6800);
   U7375 : AOI22_X1 port map( A1 => n198, A2 => n5162, B1 => n163, B2 => n5163,
                           ZN => n6798);
   U7376 : AOI22_X1 port map( A1 => n240, A2 => n5164, B1 => n160, B2 => n5165,
                           ZN => n6797);
   U7377 : NAND3_X1 port map( A1 => n6801, A2 => n6802, A3 => n6803, ZN => 
                           n12802);
   U7378 : AOI221_X1 port map( B1 => n219, B2 => n5169, C1 => n6682, C2 => 
                           MEM_IN(30), A => n6804, ZN => n6803);
   U7379 : OAI22_X1 port map( A1 => n11439, A2 => n247, B1 => n5171, B2 => n148
                           , ZN => n6804);
   U7380 : AOI22_X1 port map( A1 => n198, A2 => n5172, B1 => n163, B2 => n5173,
                           ZN => n6802);
   U7381 : AOI22_X1 port map( A1 => n240, A2 => n5174, B1 => n160, B2 => n5175,
                           ZN => n6801);
   U7382 : NAND3_X1 port map( A1 => n6805, A2 => n6806, A3 => n6807, ZN => 
                           n12801);
   U7383 : AOI221_X1 port map( B1 => n219, B2 => n5179, C1 => n6682, C2 => 
                           MEM_IN(31), A => n6808, ZN => n6807);
   U7384 : OAI22_X1 port map( A1 => n11438, A2 => n247, B1 => n5181, B2 => n148
                           , ZN => n6808);
   U7385 : INV_X1 port map( A => n6814, ZN => n6813);
   U7386 : AOI22_X1 port map( A1 => n198, A2 => n5191, B1 => n163, B2 => n5192,
                           ZN => n6806);
   U7387 : AOI22_X1 port map( A1 => n240, A2 => n5195, B1 => n160, B2 => n5196,
                           ZN => n6805);
   U7388 : INV_X1 port map( A => n6522, ZN => n6521);
   U7389 : AOI22_X1 port map( A1 => n6817, A2 => n6810, B1 => n4841, B2 => n247
                           , ZN => n6812);
   U7390 : AND3_X1 port map( A1 => n208, A2 => n247, A3 => n5773, ZN => n6810);
   U7391 : INV_X1 port map( A => n6809, ZN => n5773);
   U7392 : OAI22_X1 port map( A1 => n4786, A2 => n6818, B1 => n6819, B2 => 
                           n5204, ZN => n6684);
   U7393 : NOR2_X1 port map( A1 => n6809, A2 => n6811, ZN => n6819);
   U7394 : NAND4_X1 port map( A1 => n6676, A2 => n6678, A3 => n5925, A4 => 
                           n6820, ZN => n6809);
   U7395 : AND4_X1 port map( A1 => n6821, A2 => n6671, A3 => n5368, A4 => n6815
                           , ZN => n6818);
   U7396 : INV_X1 port map( A => n6672, ZN => n6671);
   U7397 : AOI211_X1 port map( C1 => n5522, C2 => n6527, A => n6369, B => n6522
                           , ZN => n6821);
   U7398 : NOR2_X1 port map( A1 => n5925, A2 => n4787, ZN => n6369);
   U7399 : INV_X1 port map( A => n6811, ZN => n6817);
   U7400 : NAND2_X1 port map( A1 => n6822, A2 => n6823, ZN => n6811);
   U7401 : NAND2_X1 port map( A1 => n6531, A2 => n5526, ZN => n5925);
   U7402 : NAND3_X1 port map( A1 => n6824, A2 => n6825, A3 => n6826, ZN => 
                           n12800);
   U7403 : AOI221_X1 port map( B1 => n6827, B2 => n4863, C1 => n190, C2 => 
                           MEM_IN(0), A => n6828, ZN => n6826);
   U7404 : OAI22_X1 port map( A1 => n11437, A2 => n293, B1 => n4867, B2 => n149
                           , ZN => n6828);
   U7405 : AOI22_X1 port map( A1 => n6830, A2 => n4869, B1 => n6831, B2 => 
                           n4871, ZN => n6825);
   U7406 : AOI22_X1 port map( A1 => n6832, A2 => n4873, B1 => n6833, B2 => 
                           n4875, ZN => n6824);
   U7407 : NAND3_X1 port map( A1 => n6834, A2 => n6835, A3 => n6836, ZN => 
                           n12799);
   U7408 : AOI221_X1 port map( B1 => n6827, B2 => n4879, C1 => n190, C2 => 
                           MEM_IN(1), A => n6837, ZN => n6836);
   U7409 : OAI22_X1 port map( A1 => n11436, A2 => n293, B1 => n4881, B2 => n149
                           , ZN => n6837);
   U7410 : AOI22_X1 port map( A1 => n6830, A2 => n4882, B1 => n6831, B2 => 
                           n4883, ZN => n6835);
   U7411 : AOI22_X1 port map( A1 => n6832, A2 => n4884, B1 => n6833, B2 => 
                           n4885, ZN => n6834);
   U7412 : NAND3_X1 port map( A1 => n6838, A2 => n6839, A3 => n6840, ZN => 
                           n12798);
   U7413 : AOI221_X1 port map( B1 => n6827, B2 => n4889, C1 => n190, C2 => 
                           MEM_IN(2), A => n6841, ZN => n6840);
   U7414 : OAI22_X1 port map( A1 => n11435, A2 => n293, B1 => n4891, B2 => n149
                           , ZN => n6841);
   U7415 : AOI22_X1 port map( A1 => n6830, A2 => n4892, B1 => n6831, B2 => 
                           n4893, ZN => n6839);
   U7416 : AOI22_X1 port map( A1 => n6832, A2 => n4894, B1 => n6833, B2 => 
                           n4895, ZN => n6838);
   U7417 : NAND3_X1 port map( A1 => n6842, A2 => n6843, A3 => n6844, ZN => 
                           n12797);
   U7418 : AOI221_X1 port map( B1 => n6827, B2 => n4899, C1 => n190, C2 => 
                           MEM_IN(3), A => n6845, ZN => n6844);
   U7419 : OAI22_X1 port map( A1 => n11434, A2 => n293, B1 => n4901, B2 => n149
                           , ZN => n6845);
   U7420 : AOI22_X1 port map( A1 => n6830, A2 => n4902, B1 => n6831, B2 => 
                           n4903, ZN => n6843);
   U7421 : AOI22_X1 port map( A1 => n6832, A2 => n4904, B1 => n6833, B2 => 
                           n4905, ZN => n6842);
   U7422 : NAND3_X1 port map( A1 => n6846, A2 => n6847, A3 => n6848, ZN => 
                           n12796);
   U7423 : AOI221_X1 port map( B1 => n6827, B2 => n4909, C1 => n190, C2 => 
                           MEM_IN(4), A => n6849, ZN => n6848);
   U7424 : OAI22_X1 port map( A1 => n11433, A2 => n293, B1 => n4911, B2 => n149
                           , ZN => n6849);
   U7425 : AOI22_X1 port map( A1 => n6830, A2 => n4912, B1 => n6831, B2 => 
                           n4913, ZN => n6847);
   U7426 : AOI22_X1 port map( A1 => n6832, A2 => n4914, B1 => n6833, B2 => 
                           n4915, ZN => n6846);
   U7427 : NAND3_X1 port map( A1 => n6850, A2 => n6851, A3 => n6852, ZN => 
                           n12795);
   U7428 : AOI221_X1 port map( B1 => n6827, B2 => n4919, C1 => n190, C2 => 
                           MEM_IN(5), A => n6853, ZN => n6852);
   U7429 : OAI22_X1 port map( A1 => n11432, A2 => n293, B1 => n4921, B2 => n149
                           , ZN => n6853);
   U7430 : AOI22_X1 port map( A1 => n6830, A2 => n4922, B1 => n6831, B2 => 
                           n4923, ZN => n6851);
   U7431 : AOI22_X1 port map( A1 => n6832, A2 => n4924, B1 => n6833, B2 => 
                           n4925, ZN => n6850);
   U7432 : NAND3_X1 port map( A1 => n6854, A2 => n6855, A3 => n6856, ZN => 
                           n12794);
   U7433 : AOI221_X1 port map( B1 => n6827, B2 => n4929, C1 => n190, C2 => 
                           MEM_IN(6), A => n6857, ZN => n6856);
   U7434 : OAI22_X1 port map( A1 => n11431, A2 => n293, B1 => n4931, B2 => n149
                           , ZN => n6857);
   U7435 : AOI22_X1 port map( A1 => n6830, A2 => n4932, B1 => n6831, B2 => 
                           n4933, ZN => n6855);
   U7436 : AOI22_X1 port map( A1 => n6832, A2 => n4934, B1 => n6833, B2 => 
                           n4935, ZN => n6854);
   U7437 : NAND3_X1 port map( A1 => n6858, A2 => n6859, A3 => n6860, ZN => 
                           n12793);
   U7438 : AOI221_X1 port map( B1 => n6827, B2 => n4939, C1 => n190, C2 => 
                           MEM_IN(7), A => n6861, ZN => n6860);
   U7439 : OAI22_X1 port map( A1 => n11430, A2 => n293, B1 => n4941, B2 => n149
                           , ZN => n6861);
   U7440 : AOI22_X1 port map( A1 => n6830, A2 => n4942, B1 => n6831, B2 => 
                           n4943, ZN => n6859);
   U7441 : AOI22_X1 port map( A1 => n6832, A2 => n4944, B1 => n6833, B2 => 
                           n4945, ZN => n6858);
   U7442 : NAND3_X1 port map( A1 => n6862, A2 => n6863, A3 => n6864, ZN => 
                           n12792);
   U7443 : AOI221_X1 port map( B1 => n6827, B2 => n4949, C1 => n190, C2 => 
                           MEM_IN(8), A => n6865, ZN => n6864);
   U7444 : OAI22_X1 port map( A1 => n11429, A2 => n293, B1 => n4951, B2 => n149
                           , ZN => n6865);
   U7445 : AOI22_X1 port map( A1 => n6830, A2 => n4952, B1 => n6831, B2 => 
                           n4953, ZN => n6863);
   U7446 : AOI22_X1 port map( A1 => n6832, A2 => n4954, B1 => n6833, B2 => 
                           n4955, ZN => n6862);
   U7447 : NAND3_X1 port map( A1 => n6866, A2 => n6867, A3 => n6868, ZN => 
                           n12791);
   U7448 : AOI221_X1 port map( B1 => n6827, B2 => n4959, C1 => n190, C2 => 
                           MEM_IN(9), A => n6869, ZN => n6868);
   U7449 : OAI22_X1 port map( A1 => n11428, A2 => n293, B1 => n4961, B2 => n149
                           , ZN => n6869);
   U7450 : AOI22_X1 port map( A1 => n6830, A2 => n4962, B1 => n6831, B2 => 
                           n4963, ZN => n6867);
   U7451 : AOI22_X1 port map( A1 => n6832, A2 => n4964, B1 => n6833, B2 => 
                           n4965, ZN => n6866);
   U7452 : NAND3_X1 port map( A1 => n6870, A2 => n6871, A3 => n6872, ZN => 
                           n12790);
   U7453 : AOI221_X1 port map( B1 => n6827, B2 => n4969, C1 => n190, C2 => 
                           MEM_IN(10), A => n6873, ZN => n6872);
   U7454 : OAI22_X1 port map( A1 => n11427, A2 => n293, B1 => n4971, B2 => n149
                           , ZN => n6873);
   U7455 : AOI22_X1 port map( A1 => n6830, A2 => n4972, B1 => n6831, B2 => 
                           n4973, ZN => n6871);
   U7456 : AOI22_X1 port map( A1 => n6832, A2 => n4974, B1 => n6833, B2 => 
                           n4975, ZN => n6870);
   U7457 : NAND3_X1 port map( A1 => n6874, A2 => n6875, A3 => n6876, ZN => 
                           n12789);
   U7458 : AOI221_X1 port map( B1 => n6827, B2 => n4979, C1 => n190, C2 => 
                           MEM_IN(11), A => n6877, ZN => n6876);
   U7459 : OAI22_X1 port map( A1 => n11426, A2 => n293, B1 => n4981, B2 => n149
                           , ZN => n6877);
   U7460 : AOI22_X1 port map( A1 => n6830, A2 => n4982, B1 => n6831, B2 => 
                           n4983, ZN => n6875);
   U7461 : AOI22_X1 port map( A1 => n6832, A2 => n4984, B1 => n6833, B2 => 
                           n4985, ZN => n6874);
   U7462 : NAND3_X1 port map( A1 => n6878, A2 => n6879, A3 => n6880, ZN => 
                           n12788);
   U7463 : AOI221_X1 port map( B1 => n6827, B2 => n4989, C1 => n190, C2 => 
                           MEM_IN(12), A => n6881, ZN => n6880);
   U7464 : OAI22_X1 port map( A1 => n11425, A2 => n293, B1 => n4991, B2 => n149
                           , ZN => n6881);
   U7465 : AOI22_X1 port map( A1 => n6830, A2 => n4992, B1 => n6831, B2 => 
                           n4993, ZN => n6879);
   U7466 : AOI22_X1 port map( A1 => n6832, A2 => n4994, B1 => n6833, B2 => 
                           n4995, ZN => n6878);
   U7467 : NAND3_X1 port map( A1 => n6882, A2 => n6883, A3 => n6884, ZN => 
                           n12787);
   U7468 : AOI221_X1 port map( B1 => n6827, B2 => n4999, C1 => n190, C2 => 
                           MEM_IN(13), A => n6885, ZN => n6884);
   U7469 : OAI22_X1 port map( A1 => n11424, A2 => n293, B1 => n5001, B2 => n149
                           , ZN => n6885);
   U7470 : AOI22_X1 port map( A1 => n6830, A2 => n5002, B1 => n6831, B2 => 
                           n5003, ZN => n6883);
   U7471 : AOI22_X1 port map( A1 => n6832, A2 => n5004, B1 => n6833, B2 => 
                           n5005, ZN => n6882);
   U7472 : NAND3_X1 port map( A1 => n6886, A2 => n6887, A3 => n6888, ZN => 
                           n12786);
   U7473 : AOI221_X1 port map( B1 => n6827, B2 => n5009, C1 => n190, C2 => 
                           MEM_IN(14), A => n6889, ZN => n6888);
   U7474 : OAI22_X1 port map( A1 => n11423, A2 => n293, B1 => n5011, B2 => n149
                           , ZN => n6889);
   U7475 : AOI22_X1 port map( A1 => n6830, A2 => n5012, B1 => n6831, B2 => 
                           n5013, ZN => n6887);
   U7476 : AOI22_X1 port map( A1 => n6832, A2 => n5014, B1 => n6833, B2 => 
                           n5015, ZN => n6886);
   U7477 : NAND3_X1 port map( A1 => n6890, A2 => n6891, A3 => n6892, ZN => 
                           n12785);
   U7478 : AOI221_X1 port map( B1 => n6827, B2 => n5019, C1 => n190, C2 => 
                           MEM_IN(15), A => n6893, ZN => n6892);
   U7479 : OAI22_X1 port map( A1 => n11422, A2 => n293, B1 => n5021, B2 => n149
                           , ZN => n6893);
   U7480 : AOI22_X1 port map( A1 => n6830, A2 => n5022, B1 => n6831, B2 => 
                           n5023, ZN => n6891);
   U7481 : AOI22_X1 port map( A1 => n6832, A2 => n5024, B1 => n6833, B2 => 
                           n5025, ZN => n6890);
   U7482 : NAND3_X1 port map( A1 => n6894, A2 => n6895, A3 => n6896, ZN => 
                           n12784);
   U7483 : AOI221_X1 port map( B1 => n6827, B2 => n5029, C1 => n190, C2 => 
                           MEM_IN(16), A => n6897, ZN => n6896);
   U7484 : OAI22_X1 port map( A1 => n11421, A2 => n293, B1 => n5031, B2 => n149
                           , ZN => n6897);
   U7485 : AOI22_X1 port map( A1 => n6830, A2 => n5032, B1 => n6831, B2 => 
                           n5033, ZN => n6895);
   U7486 : AOI22_X1 port map( A1 => n6832, A2 => n5034, B1 => n6833, B2 => 
                           n5035, ZN => n6894);
   U7487 : NAND3_X1 port map( A1 => n6898, A2 => n6899, A3 => n6900, ZN => 
                           n12783);
   U7488 : AOI221_X1 port map( B1 => n6827, B2 => n5039, C1 => n190, C2 => 
                           MEM_IN(17), A => n6901, ZN => n6900);
   U7489 : OAI22_X1 port map( A1 => n11420, A2 => n293, B1 => n5041, B2 => n149
                           , ZN => n6901);
   U7490 : AOI22_X1 port map( A1 => n6830, A2 => n5042, B1 => n6831, B2 => 
                           n5043, ZN => n6899);
   U7491 : AOI22_X1 port map( A1 => n6832, A2 => n5044, B1 => n6833, B2 => 
                           n5045, ZN => n6898);
   U7492 : NAND3_X1 port map( A1 => n6902, A2 => n6903, A3 => n6904, ZN => 
                           n12782);
   U7493 : AOI221_X1 port map( B1 => n6827, B2 => n5049, C1 => n190, C2 => 
                           MEM_IN(18), A => n6905, ZN => n6904);
   U7494 : OAI22_X1 port map( A1 => n11419, A2 => n293, B1 => n5051, B2 => n149
                           , ZN => n6905);
   U7495 : AOI22_X1 port map( A1 => n6830, A2 => n5052, B1 => n6831, B2 => 
                           n5053, ZN => n6903);
   U7496 : AOI22_X1 port map( A1 => n6832, A2 => n5054, B1 => n6833, B2 => 
                           n5055, ZN => n6902);
   U7497 : NAND3_X1 port map( A1 => n6906, A2 => n6907, A3 => n6908, ZN => 
                           n12781);
   U7498 : AOI221_X1 port map( B1 => n6827, B2 => n5059, C1 => n190, C2 => 
                           MEM_IN(19), A => n6909, ZN => n6908);
   U7499 : OAI22_X1 port map( A1 => n11418, A2 => n293, B1 => n5061, B2 => n149
                           , ZN => n6909);
   U7500 : AOI22_X1 port map( A1 => n6830, A2 => n5062, B1 => n6831, B2 => 
                           n5063, ZN => n6907);
   U7501 : AOI22_X1 port map( A1 => n6832, A2 => n5064, B1 => n6833, B2 => 
                           n5065, ZN => n6906);
   U7502 : NAND3_X1 port map( A1 => n6910, A2 => n6911, A3 => n6912, ZN => 
                           n12780);
   U7503 : AOI221_X1 port map( B1 => n6827, B2 => n5069, C1 => n190, C2 => 
                           MEM_IN(20), A => n6913, ZN => n6912);
   U7504 : OAI22_X1 port map( A1 => n11417, A2 => n293, B1 => n5071, B2 => n149
                           , ZN => n6913);
   U7505 : AOI22_X1 port map( A1 => n6830, A2 => n5072, B1 => n6831, B2 => 
                           n5073, ZN => n6911);
   U7506 : AOI22_X1 port map( A1 => n6832, A2 => n5074, B1 => n6833, B2 => 
                           n5075, ZN => n6910);
   U7507 : NAND3_X1 port map( A1 => n6914, A2 => n6915, A3 => n6916, ZN => 
                           n12779);
   U7508 : AOI221_X1 port map( B1 => n6827, B2 => n5079, C1 => n190, C2 => 
                           MEM_IN(21), A => n6917, ZN => n6916);
   U7509 : OAI22_X1 port map( A1 => n11416, A2 => n293, B1 => n5081, B2 => n149
                           , ZN => n6917);
   U7510 : AOI22_X1 port map( A1 => n6830, A2 => n5082, B1 => n6831, B2 => 
                           n5083, ZN => n6915);
   U7511 : AOI22_X1 port map( A1 => n6832, A2 => n5084, B1 => n6833, B2 => 
                           n5085, ZN => n6914);
   U7512 : NAND3_X1 port map( A1 => n6918, A2 => n6919, A3 => n6920, ZN => 
                           n12778);
   U7513 : AOI221_X1 port map( B1 => n6827, B2 => n5089, C1 => n190, C2 => 
                           MEM_IN(22), A => n6921, ZN => n6920);
   U7514 : OAI22_X1 port map( A1 => n11415, A2 => n293, B1 => n5091, B2 => n149
                           , ZN => n6921);
   U7515 : AOI22_X1 port map( A1 => n6830, A2 => n5092, B1 => n6831, B2 => 
                           n5093, ZN => n6919);
   U7516 : AOI22_X1 port map( A1 => n6832, A2 => n5094, B1 => n6833, B2 => 
                           n5095, ZN => n6918);
   U7517 : NAND3_X1 port map( A1 => n6922, A2 => n6923, A3 => n6924, ZN => 
                           n12777);
   U7518 : AOI221_X1 port map( B1 => n6827, B2 => n5099, C1 => n190, C2 => 
                           MEM_IN(23), A => n6925, ZN => n6924);
   U7519 : OAI22_X1 port map( A1 => n11414, A2 => n293, B1 => n5101, B2 => n149
                           , ZN => n6925);
   U7520 : AOI22_X1 port map( A1 => n6830, A2 => n5102, B1 => n6831, B2 => 
                           n5103, ZN => n6923);
   U7521 : AOI22_X1 port map( A1 => n6832, A2 => n5104, B1 => n6833, B2 => 
                           n5105, ZN => n6922);
   U7522 : NAND3_X1 port map( A1 => n6926, A2 => n6927, A3 => n6928, ZN => 
                           n12776);
   U7523 : AOI221_X1 port map( B1 => n6827, B2 => n5109, C1 => n190, C2 => 
                           MEM_IN(24), A => n6929, ZN => n6928);
   U7524 : OAI22_X1 port map( A1 => n11413, A2 => n293, B1 => n5111, B2 => n149
                           , ZN => n6929);
   U7525 : AOI22_X1 port map( A1 => n6830, A2 => n5112, B1 => n6831, B2 => 
                           n5113, ZN => n6927);
   U7526 : AOI22_X1 port map( A1 => n6832, A2 => n5114, B1 => n6833, B2 => 
                           n5115, ZN => n6926);
   U7527 : NAND3_X1 port map( A1 => n6930, A2 => n6931, A3 => n6932, ZN => 
                           n12775);
   U7528 : AOI221_X1 port map( B1 => n6827, B2 => n5119, C1 => n190, C2 => 
                           MEM_IN(25), A => n6933, ZN => n6932);
   U7529 : OAI22_X1 port map( A1 => n11412, A2 => n293, B1 => n5121, B2 => n149
                           , ZN => n6933);
   U7530 : AOI22_X1 port map( A1 => n6830, A2 => n5122, B1 => n6831, B2 => 
                           n5123, ZN => n6931);
   U7531 : AOI22_X1 port map( A1 => n6832, A2 => n5124, B1 => n6833, B2 => 
                           n5125, ZN => n6930);
   U7532 : NAND3_X1 port map( A1 => n6934, A2 => n6935, A3 => n6936, ZN => 
                           n12774);
   U7533 : AOI221_X1 port map( B1 => n6827, B2 => n5129, C1 => n190, C2 => 
                           MEM_IN(26), A => n6937, ZN => n6936);
   U7534 : OAI22_X1 port map( A1 => n11411, A2 => n293, B1 => n5131, B2 => n149
                           , ZN => n6937);
   U7535 : AOI22_X1 port map( A1 => n6830, A2 => n5132, B1 => n6831, B2 => 
                           n5133, ZN => n6935);
   U7536 : AOI22_X1 port map( A1 => n6832, A2 => n5134, B1 => n6833, B2 => 
                           n5135, ZN => n6934);
   U7537 : NAND3_X1 port map( A1 => n6938, A2 => n6939, A3 => n6940, ZN => 
                           n12773);
   U7538 : AOI221_X1 port map( B1 => n6827, B2 => n5139, C1 => n190, C2 => 
                           MEM_IN(27), A => n6941, ZN => n6940);
   U7539 : OAI22_X1 port map( A1 => n11410, A2 => n293, B1 => n5141, B2 => n149
                           , ZN => n6941);
   U7540 : AOI22_X1 port map( A1 => n6830, A2 => n5142, B1 => n6831, B2 => 
                           n5143, ZN => n6939);
   U7541 : AOI22_X1 port map( A1 => n6832, A2 => n5144, B1 => n6833, B2 => 
                           n5145, ZN => n6938);
   U7542 : NAND3_X1 port map( A1 => n6942, A2 => n6943, A3 => n6944, ZN => 
                           n12772);
   U7543 : AOI221_X1 port map( B1 => n6827, B2 => n5149, C1 => n190, C2 => 
                           MEM_IN(28), A => n6945, ZN => n6944);
   U7544 : OAI22_X1 port map( A1 => n11409, A2 => n293, B1 => n5151, B2 => n149
                           , ZN => n6945);
   U7545 : AOI22_X1 port map( A1 => n6830, A2 => n5152, B1 => n6831, B2 => 
                           n5153, ZN => n6943);
   U7546 : AOI22_X1 port map( A1 => n6832, A2 => n5154, B1 => n6833, B2 => 
                           n5155, ZN => n6942);
   U7547 : NAND3_X1 port map( A1 => n6946, A2 => n6947, A3 => n6948, ZN => 
                           n12771);
   U7548 : AOI221_X1 port map( B1 => n6827, B2 => n5159, C1 => n190, C2 => 
                           MEM_IN(29), A => n6949, ZN => n6948);
   U7549 : OAI22_X1 port map( A1 => n11408, A2 => n293, B1 => n5161, B2 => n149
                           , ZN => n6949);
   U7550 : AOI22_X1 port map( A1 => n6830, A2 => n5162, B1 => n6831, B2 => 
                           n5163, ZN => n6947);
   U7551 : AOI22_X1 port map( A1 => n6832, A2 => n5164, B1 => n6833, B2 => 
                           n5165, ZN => n6946);
   U7552 : NAND3_X1 port map( A1 => n6950, A2 => n6951, A3 => n6952, ZN => 
                           n12770);
   U7553 : AOI221_X1 port map( B1 => n6827, B2 => n5169, C1 => n190, C2 => 
                           MEM_IN(30), A => n6953, ZN => n6952);
   U7554 : OAI22_X1 port map( A1 => n11407, A2 => n293, B1 => n5171, B2 => n149
                           , ZN => n6953);
   U7555 : AOI22_X1 port map( A1 => n6830, A2 => n5172, B1 => n6831, B2 => 
                           n5173, ZN => n6951);
   U7556 : AOI22_X1 port map( A1 => n6832, A2 => n5174, B1 => n6833, B2 => 
                           n5175, ZN => n6950);
   U7557 : NAND3_X1 port map( A1 => n6954, A2 => n6955, A3 => n6956, ZN => 
                           n12769);
   U7558 : AOI221_X1 port map( B1 => n6827, B2 => n5179, C1 => n190, C2 => 
                           MEM_IN(31), A => n6957, ZN => n6956);
   U7559 : OAI22_X1 port map( A1 => n11406, A2 => n293, B1 => n5181, B2 => n149
                           , ZN => n6957);
   U7560 : NAND2_X1 port map( A1 => n5206, A2 => n6816, ZN => n6814);
   U7561 : NAND3_X1 port map( A1 => n5206, A2 => n6820, A3 => n6526, ZN => 
                           n6816);
   U7562 : AOI22_X1 port map( A1 => n6830, A2 => n5191, B1 => n6831, B2 => 
                           n5192, ZN => n6955);
   U7563 : AOI22_X1 port map( A1 => n6832, A2 => n5195, B1 => n6833, B2 => 
                           n5196, ZN => n6954);
   U7564 : OAI22_X1 port map( A1 => n6965, A2 => n6959, B1 => n208, B2 => n292,
                           ZN => n6962);
   U7565 : NAND3_X1 port map( A1 => n208, A2 => n293, A3 => n5924, ZN => n6959)
                           ;
   U7566 : OAI22_X1 port map( A1 => n4786, A2 => n6966, B1 => n6967, B2 => 
                           n5204, ZN => n6829);
   U7567 : NOR2_X1 port map( A1 => n6958, A2 => n6965, ZN => n6967);
   U7568 : INV_X1 port map( A => n5924, ZN => n6958);
   U7569 : NOR3_X1 port map( A1 => n6968, A2 => n6078, A3 => n6969, ZN => n5924
                           );
   U7570 : INV_X1 port map( A => n6820, ZN => n6078);
   U7571 : NOR3_X1 port map( A1 => n6970, A2 => RESET, A3 => n6522, ZN => n6966
                           );
   U7572 : OAI22_X1 port map( A1 => n5771, A2 => n6971, B1 => n6676, B2 => 
                           n4787, ZN => n6970);
   U7573 : INV_X1 port map( A => n6960, ZN => n6965);
   U7574 : NOR2_X1 port map( A1 => n6972, A2 => n6973, ZN => n6960);
   U7575 : NOR2_X1 port map( A1 => n6820, A2 => n4787, ZN => n6522);
   U7576 : NAND2_X1 port map( A1 => n6531, A2 => n5775, ZN => n6820);
   U7577 : NAND3_X1 port map( A1 => n6974, A2 => n6975, A3 => n6976, ZN => 
                           n12768);
   U7578 : AOI221_X1 port map( B1 => n6977, B2 => n4863, C1 => n6978, C2 => 
                           MEM_IN(0), A => n6979, ZN => n6976);
   U7579 : OAI22_X1 port map( A1 => n11405, A2 => n216, B1 => n4867, B2 => n146
                           , ZN => n6979);
   U7580 : AOI22_X1 port map( A1 => n6981, A2 => n4869, B1 => n6982, B2 => 
                           n4871, ZN => n6975);
   U7581 : AOI22_X1 port map( A1 => n6983, A2 => n4873, B1 => n6984, B2 => 
                           n4875, ZN => n6974);
   U7582 : NAND3_X1 port map( A1 => n6985, A2 => n6986, A3 => n6987, ZN => 
                           n12767);
   U7583 : AOI221_X1 port map( B1 => n6977, B2 => n4879, C1 => n6978, C2 => 
                           MEM_IN(1), A => n6988, ZN => n6987);
   U7584 : OAI22_X1 port map( A1 => n11404, A2 => n216, B1 => n4881, B2 => n146
                           , ZN => n6988);
   U7585 : AOI22_X1 port map( A1 => n6981, A2 => n4882, B1 => n6982, B2 => 
                           n4883, ZN => n6986);
   U7586 : AOI22_X1 port map( A1 => n6983, A2 => n4884, B1 => n6984, B2 => 
                           n4885, ZN => n6985);
   U7587 : NAND3_X1 port map( A1 => n6989, A2 => n6990, A3 => n6991, ZN => 
                           n12766);
   U7588 : AOI221_X1 port map( B1 => n6977, B2 => n4889, C1 => n6978, C2 => 
                           MEM_IN(2), A => n6992, ZN => n6991);
   U7589 : OAI22_X1 port map( A1 => n11403, A2 => n216, B1 => n4891, B2 => n146
                           , ZN => n6992);
   U7590 : AOI22_X1 port map( A1 => n6981, A2 => n4892, B1 => n6982, B2 => 
                           n4893, ZN => n6990);
   U7591 : AOI22_X1 port map( A1 => n6983, A2 => n4894, B1 => n6984, B2 => 
                           n4895, ZN => n6989);
   U7592 : NAND3_X1 port map( A1 => n6993, A2 => n6994, A3 => n6995, ZN => 
                           n12765);
   U7593 : AOI221_X1 port map( B1 => n6977, B2 => n4899, C1 => n6978, C2 => 
                           MEM_IN(3), A => n6996, ZN => n6995);
   U7594 : OAI22_X1 port map( A1 => n11402, A2 => n216, B1 => n4901, B2 => n146
                           , ZN => n6996);
   U7595 : AOI22_X1 port map( A1 => n6981, A2 => n4902, B1 => n6982, B2 => 
                           n4903, ZN => n6994);
   U7596 : AOI22_X1 port map( A1 => n6983, A2 => n4904, B1 => n6984, B2 => 
                           n4905, ZN => n6993);
   U7597 : NAND3_X1 port map( A1 => n6997, A2 => n6998, A3 => n6999, ZN => 
                           n12764);
   U7598 : AOI221_X1 port map( B1 => n6977, B2 => n4909, C1 => n6978, C2 => 
                           MEM_IN(4), A => n7000, ZN => n6999);
   U7599 : OAI22_X1 port map( A1 => n11401, A2 => n216, B1 => n4911, B2 => n146
                           , ZN => n7000);
   U7600 : AOI22_X1 port map( A1 => n6981, A2 => n4912, B1 => n6982, B2 => 
                           n4913, ZN => n6998);
   U7601 : AOI22_X1 port map( A1 => n6983, A2 => n4914, B1 => n6984, B2 => 
                           n4915, ZN => n6997);
   U7602 : NAND3_X1 port map( A1 => n7001, A2 => n7002, A3 => n7003, ZN => 
                           n12763);
   U7603 : AOI221_X1 port map( B1 => n6977, B2 => n4919, C1 => n6978, C2 => 
                           MEM_IN(5), A => n7004, ZN => n7003);
   U7604 : OAI22_X1 port map( A1 => n11400, A2 => n216, B1 => n4921, B2 => n146
                           , ZN => n7004);
   U7605 : AOI22_X1 port map( A1 => n6981, A2 => n4922, B1 => n6982, B2 => 
                           n4923, ZN => n7002);
   U7606 : AOI22_X1 port map( A1 => n6983, A2 => n4924, B1 => n6984, B2 => 
                           n4925, ZN => n7001);
   U7607 : NAND3_X1 port map( A1 => n7005, A2 => n7006, A3 => n7007, ZN => 
                           n12762);
   U7608 : AOI221_X1 port map( B1 => n6977, B2 => n4929, C1 => n6978, C2 => 
                           MEM_IN(6), A => n7008, ZN => n7007);
   U7609 : OAI22_X1 port map( A1 => n11399, A2 => n216, B1 => n4931, B2 => n146
                           , ZN => n7008);
   U7610 : AOI22_X1 port map( A1 => n6981, A2 => n4932, B1 => n6982, B2 => 
                           n4933, ZN => n7006);
   U7611 : AOI22_X1 port map( A1 => n6983, A2 => n4934, B1 => n6984, B2 => 
                           n4935, ZN => n7005);
   U7612 : NAND3_X1 port map( A1 => n7009, A2 => n7010, A3 => n7011, ZN => 
                           n12761);
   U7613 : AOI221_X1 port map( B1 => n6977, B2 => n4939, C1 => n6978, C2 => 
                           MEM_IN(7), A => n7012, ZN => n7011);
   U7614 : OAI22_X1 port map( A1 => n11398, A2 => n216, B1 => n4941, B2 => n146
                           , ZN => n7012);
   U7615 : AOI22_X1 port map( A1 => n6981, A2 => n4942, B1 => n6982, B2 => 
                           n4943, ZN => n7010);
   U7616 : AOI22_X1 port map( A1 => n6983, A2 => n4944, B1 => n6984, B2 => 
                           n4945, ZN => n7009);
   U7617 : NAND3_X1 port map( A1 => n7013, A2 => n7014, A3 => n7015, ZN => 
                           n12760);
   U7618 : AOI221_X1 port map( B1 => n6977, B2 => n4949, C1 => n6978, C2 => 
                           MEM_IN(8), A => n7016, ZN => n7015);
   U7619 : OAI22_X1 port map( A1 => n11397, A2 => n216, B1 => n4951, B2 => n146
                           , ZN => n7016);
   U7620 : AOI22_X1 port map( A1 => n6981, A2 => n4952, B1 => n6982, B2 => 
                           n4953, ZN => n7014);
   U7621 : AOI22_X1 port map( A1 => n6983, A2 => n4954, B1 => n6984, B2 => 
                           n4955, ZN => n7013);
   U7622 : NAND3_X1 port map( A1 => n7017, A2 => n7018, A3 => n7019, ZN => 
                           n12759);
   U7623 : AOI221_X1 port map( B1 => n6977, B2 => n4959, C1 => n6978, C2 => 
                           MEM_IN(9), A => n7020, ZN => n7019);
   U7624 : OAI22_X1 port map( A1 => n11396, A2 => n216, B1 => n4961, B2 => n146
                           , ZN => n7020);
   U7625 : AOI22_X1 port map( A1 => n6981, A2 => n4962, B1 => n6982, B2 => 
                           n4963, ZN => n7018);
   U7626 : AOI22_X1 port map( A1 => n6983, A2 => n4964, B1 => n6984, B2 => 
                           n4965, ZN => n7017);
   U7627 : NAND3_X1 port map( A1 => n7021, A2 => n7022, A3 => n7023, ZN => 
                           n12758);
   U7628 : AOI221_X1 port map( B1 => n6977, B2 => n4969, C1 => n6978, C2 => 
                           MEM_IN(10), A => n7024, ZN => n7023);
   U7629 : OAI22_X1 port map( A1 => n11395, A2 => n216, B1 => n4971, B2 => n146
                           , ZN => n7024);
   U7630 : AOI22_X1 port map( A1 => n6981, A2 => n4972, B1 => n6982, B2 => 
                           n4973, ZN => n7022);
   U7631 : AOI22_X1 port map( A1 => n6983, A2 => n4974, B1 => n6984, B2 => 
                           n4975, ZN => n7021);
   U7632 : NAND3_X1 port map( A1 => n7025, A2 => n7026, A3 => n7027, ZN => 
                           n12757);
   U7633 : AOI221_X1 port map( B1 => n6977, B2 => n4979, C1 => n6978, C2 => 
                           MEM_IN(11), A => n7028, ZN => n7027);
   U7634 : OAI22_X1 port map( A1 => n11394, A2 => n216, B1 => n4981, B2 => n146
                           , ZN => n7028);
   U7635 : AOI22_X1 port map( A1 => n6981, A2 => n4982, B1 => n6982, B2 => 
                           n4983, ZN => n7026);
   U7636 : AOI22_X1 port map( A1 => n6983, A2 => n4984, B1 => n6984, B2 => 
                           n4985, ZN => n7025);
   U7637 : NAND3_X1 port map( A1 => n7029, A2 => n7030, A3 => n7031, ZN => 
                           n12756);
   U7638 : AOI221_X1 port map( B1 => n6977, B2 => n4989, C1 => n6978, C2 => 
                           MEM_IN(12), A => n7032, ZN => n7031);
   U7639 : OAI22_X1 port map( A1 => n11393, A2 => n216, B1 => n4991, B2 => n146
                           , ZN => n7032);
   U7640 : AOI22_X1 port map( A1 => n6981, A2 => n4992, B1 => n6982, B2 => 
                           n4993, ZN => n7030);
   U7641 : AOI22_X1 port map( A1 => n6983, A2 => n4994, B1 => n6984, B2 => 
                           n4995, ZN => n7029);
   U7642 : NAND3_X1 port map( A1 => n7033, A2 => n7034, A3 => n7035, ZN => 
                           n12755);
   U7643 : AOI221_X1 port map( B1 => n6977, B2 => n4999, C1 => n6978, C2 => 
                           MEM_IN(13), A => n7036, ZN => n7035);
   U7644 : OAI22_X1 port map( A1 => n11392, A2 => n216, B1 => n5001, B2 => n146
                           , ZN => n7036);
   U7645 : AOI22_X1 port map( A1 => n6981, A2 => n5002, B1 => n6982, B2 => 
                           n5003, ZN => n7034);
   U7646 : AOI22_X1 port map( A1 => n6983, A2 => n5004, B1 => n6984, B2 => 
                           n5005, ZN => n7033);
   U7647 : NAND3_X1 port map( A1 => n7037, A2 => n7038, A3 => n7039, ZN => 
                           n12754);
   U7648 : AOI221_X1 port map( B1 => n6977, B2 => n5009, C1 => n6978, C2 => 
                           MEM_IN(14), A => n7040, ZN => n7039);
   U7649 : OAI22_X1 port map( A1 => n11391, A2 => n216, B1 => n5011, B2 => n146
                           , ZN => n7040);
   U7650 : AOI22_X1 port map( A1 => n6981, A2 => n5012, B1 => n6982, B2 => 
                           n5013, ZN => n7038);
   U7651 : AOI22_X1 port map( A1 => n6983, A2 => n5014, B1 => n6984, B2 => 
                           n5015, ZN => n7037);
   U7652 : NAND3_X1 port map( A1 => n7041, A2 => n7042, A3 => n7043, ZN => 
                           n12753);
   U7653 : AOI221_X1 port map( B1 => n6977, B2 => n5019, C1 => n6978, C2 => 
                           MEM_IN(15), A => n7044, ZN => n7043);
   U7654 : OAI22_X1 port map( A1 => n11390, A2 => n216, B1 => n5021, B2 => n146
                           , ZN => n7044);
   U7655 : AOI22_X1 port map( A1 => n6981, A2 => n5022, B1 => n6982, B2 => 
                           n5023, ZN => n7042);
   U7656 : AOI22_X1 port map( A1 => n6983, A2 => n5024, B1 => n6984, B2 => 
                           n5025, ZN => n7041);
   U7657 : NAND3_X1 port map( A1 => n7045, A2 => n7046, A3 => n7047, ZN => 
                           n12752);
   U7658 : AOI221_X1 port map( B1 => n6977, B2 => n5029, C1 => n6978, C2 => 
                           MEM_IN(16), A => n7048, ZN => n7047);
   U7659 : OAI22_X1 port map( A1 => n11389, A2 => n216, B1 => n5031, B2 => n146
                           , ZN => n7048);
   U7660 : AOI22_X1 port map( A1 => n6981, A2 => n5032, B1 => n6982, B2 => 
                           n5033, ZN => n7046);
   U7661 : AOI22_X1 port map( A1 => n6983, A2 => n5034, B1 => n6984, B2 => 
                           n5035, ZN => n7045);
   U7662 : NAND3_X1 port map( A1 => n7049, A2 => n7050, A3 => n7051, ZN => 
                           n12751);
   U7663 : AOI221_X1 port map( B1 => n6977, B2 => n5039, C1 => n6978, C2 => 
                           MEM_IN(17), A => n7052, ZN => n7051);
   U7664 : OAI22_X1 port map( A1 => n11388, A2 => n216, B1 => n5041, B2 => n146
                           , ZN => n7052);
   U7665 : AOI22_X1 port map( A1 => n6981, A2 => n5042, B1 => n6982, B2 => 
                           n5043, ZN => n7050);
   U7666 : AOI22_X1 port map( A1 => n6983, A2 => n5044, B1 => n6984, B2 => 
                           n5045, ZN => n7049);
   U7667 : NAND3_X1 port map( A1 => n7053, A2 => n7054, A3 => n7055, ZN => 
                           n12750);
   U7668 : AOI221_X1 port map( B1 => n6977, B2 => n5049, C1 => n6978, C2 => 
                           MEM_IN(18), A => n7056, ZN => n7055);
   U7669 : OAI22_X1 port map( A1 => n11387, A2 => n216, B1 => n5051, B2 => n146
                           , ZN => n7056);
   U7670 : AOI22_X1 port map( A1 => n6981, A2 => n5052, B1 => n6982, B2 => 
                           n5053, ZN => n7054);
   U7671 : AOI22_X1 port map( A1 => n6983, A2 => n5054, B1 => n6984, B2 => 
                           n5055, ZN => n7053);
   U7672 : NAND3_X1 port map( A1 => n7057, A2 => n7058, A3 => n7059, ZN => 
                           n12749);
   U7673 : AOI221_X1 port map( B1 => n6977, B2 => n5059, C1 => n6978, C2 => 
                           MEM_IN(19), A => n7060, ZN => n7059);
   U7674 : OAI22_X1 port map( A1 => n11386, A2 => n216, B1 => n5061, B2 => n146
                           , ZN => n7060);
   U7675 : AOI22_X1 port map( A1 => n6981, A2 => n5062, B1 => n6982, B2 => 
                           n5063, ZN => n7058);
   U7676 : AOI22_X1 port map( A1 => n6983, A2 => n5064, B1 => n6984, B2 => 
                           n5065, ZN => n7057);
   U7677 : NAND3_X1 port map( A1 => n7061, A2 => n7062, A3 => n7063, ZN => 
                           n12748);
   U7678 : AOI221_X1 port map( B1 => n6977, B2 => n5069, C1 => n6978, C2 => 
                           MEM_IN(20), A => n7064, ZN => n7063);
   U7679 : OAI22_X1 port map( A1 => n11385, A2 => n216, B1 => n5071, B2 => n146
                           , ZN => n7064);
   U7680 : AOI22_X1 port map( A1 => n6981, A2 => n5072, B1 => n6982, B2 => 
                           n5073, ZN => n7062);
   U7681 : AOI22_X1 port map( A1 => n6983, A2 => n5074, B1 => n6984, B2 => 
                           n5075, ZN => n7061);
   U7682 : NAND3_X1 port map( A1 => n7065, A2 => n7066, A3 => n7067, ZN => 
                           n12747);
   U7683 : AOI221_X1 port map( B1 => n6977, B2 => n5079, C1 => n6978, C2 => 
                           MEM_IN(21), A => n7068, ZN => n7067);
   U7684 : OAI22_X1 port map( A1 => n11384, A2 => n216, B1 => n5081, B2 => n146
                           , ZN => n7068);
   U7685 : AOI22_X1 port map( A1 => n6981, A2 => n5082, B1 => n6982, B2 => 
                           n5083, ZN => n7066);
   U7686 : AOI22_X1 port map( A1 => n6983, A2 => n5084, B1 => n6984, B2 => 
                           n5085, ZN => n7065);
   U7687 : NAND3_X1 port map( A1 => n7069, A2 => n7070, A3 => n7071, ZN => 
                           n12746);
   U7688 : AOI221_X1 port map( B1 => n6977, B2 => n5089, C1 => n6978, C2 => 
                           MEM_IN(22), A => n7072, ZN => n7071);
   U7689 : OAI22_X1 port map( A1 => n11383, A2 => n216, B1 => n5091, B2 => n146
                           , ZN => n7072);
   U7690 : AOI22_X1 port map( A1 => n6981, A2 => n5092, B1 => n6982, B2 => 
                           n5093, ZN => n7070);
   U7691 : AOI22_X1 port map( A1 => n6983, A2 => n5094, B1 => n6984, B2 => 
                           n5095, ZN => n7069);
   U7692 : NAND3_X1 port map( A1 => n7073, A2 => n7074, A3 => n7075, ZN => 
                           n12745);
   U7693 : AOI221_X1 port map( B1 => n6977, B2 => n5099, C1 => n6978, C2 => 
                           MEM_IN(23), A => n7076, ZN => n7075);
   U7694 : OAI22_X1 port map( A1 => n11382, A2 => n216, B1 => n5101, B2 => n146
                           , ZN => n7076);
   U7695 : AOI22_X1 port map( A1 => n6981, A2 => n5102, B1 => n6982, B2 => 
                           n5103, ZN => n7074);
   U7696 : AOI22_X1 port map( A1 => n6983, A2 => n5104, B1 => n6984, B2 => 
                           n5105, ZN => n7073);
   U7697 : NAND3_X1 port map( A1 => n7077, A2 => n7078, A3 => n7079, ZN => 
                           n12744);
   U7698 : AOI221_X1 port map( B1 => n6977, B2 => n5109, C1 => n6978, C2 => 
                           MEM_IN(24), A => n7080, ZN => n7079);
   U7699 : OAI22_X1 port map( A1 => n11381, A2 => n216, B1 => n5111, B2 => n146
                           , ZN => n7080);
   U7700 : AOI22_X1 port map( A1 => n6981, A2 => n5112, B1 => n6982, B2 => 
                           n5113, ZN => n7078);
   U7701 : AOI22_X1 port map( A1 => n6983, A2 => n5114, B1 => n6984, B2 => 
                           n5115, ZN => n7077);
   U7702 : NAND3_X1 port map( A1 => n7081, A2 => n7082, A3 => n7083, ZN => 
                           n12743);
   U7703 : AOI221_X1 port map( B1 => n6977, B2 => n5119, C1 => n6978, C2 => 
                           MEM_IN(25), A => n7084, ZN => n7083);
   U7704 : OAI22_X1 port map( A1 => n11380, A2 => n216, B1 => n5121, B2 => n146
                           , ZN => n7084);
   U7705 : AOI22_X1 port map( A1 => n6981, A2 => n5122, B1 => n6982, B2 => 
                           n5123, ZN => n7082);
   U7706 : AOI22_X1 port map( A1 => n6983, A2 => n5124, B1 => n6984, B2 => 
                           n5125, ZN => n7081);
   U7707 : NAND3_X1 port map( A1 => n7085, A2 => n7086, A3 => n7087, ZN => 
                           n12742);
   U7708 : AOI221_X1 port map( B1 => n6977, B2 => n5129, C1 => n6978, C2 => 
                           MEM_IN(26), A => n7088, ZN => n7087);
   U7709 : OAI22_X1 port map( A1 => n11379, A2 => n216, B1 => n5131, B2 => n146
                           , ZN => n7088);
   U7710 : AOI22_X1 port map( A1 => n6981, A2 => n5132, B1 => n6982, B2 => 
                           n5133, ZN => n7086);
   U7711 : AOI22_X1 port map( A1 => n6983, A2 => n5134, B1 => n6984, B2 => 
                           n5135, ZN => n7085);
   U7712 : NAND3_X1 port map( A1 => n7089, A2 => n7090, A3 => n7091, ZN => 
                           n12741);
   U7713 : AOI221_X1 port map( B1 => n6977, B2 => n5139, C1 => n6978, C2 => 
                           MEM_IN(27), A => n7092, ZN => n7091);
   U7714 : OAI22_X1 port map( A1 => n11378, A2 => n216, B1 => n5141, B2 => n146
                           , ZN => n7092);
   U7715 : AOI22_X1 port map( A1 => n6981, A2 => n5142, B1 => n6982, B2 => 
                           n5143, ZN => n7090);
   U7716 : AOI22_X1 port map( A1 => n6983, A2 => n5144, B1 => n6984, B2 => 
                           n5145, ZN => n7089);
   U7717 : NAND3_X1 port map( A1 => n7093, A2 => n7094, A3 => n7095, ZN => 
                           n12740);
   U7718 : AOI221_X1 port map( B1 => n6977, B2 => n5149, C1 => n6978, C2 => 
                           MEM_IN(28), A => n7096, ZN => n7095);
   U7719 : OAI22_X1 port map( A1 => n11377, A2 => n216, B1 => n5151, B2 => n146
                           , ZN => n7096);
   U7720 : AOI22_X1 port map( A1 => n6981, A2 => n5152, B1 => n6982, B2 => 
                           n5153, ZN => n7094);
   U7721 : AOI22_X1 port map( A1 => n6983, A2 => n5154, B1 => n6984, B2 => 
                           n5155, ZN => n7093);
   U7722 : NAND3_X1 port map( A1 => n7097, A2 => n7098, A3 => n7099, ZN => 
                           n12739);
   U7723 : AOI221_X1 port map( B1 => n6977, B2 => n5159, C1 => n6978, C2 => 
                           MEM_IN(29), A => n7100, ZN => n7099);
   U7724 : OAI22_X1 port map( A1 => n11376, A2 => n216, B1 => n5161, B2 => n146
                           , ZN => n7100);
   U7725 : AOI22_X1 port map( A1 => n6981, A2 => n5162, B1 => n6982, B2 => 
                           n5163, ZN => n7098);
   U7726 : AOI22_X1 port map( A1 => n6983, A2 => n5164, B1 => n6984, B2 => 
                           n5165, ZN => n7097);
   U7727 : NAND3_X1 port map( A1 => n7101, A2 => n7102, A3 => n7103, ZN => 
                           n12738);
   U7728 : AOI221_X1 port map( B1 => n6977, B2 => n5169, C1 => n6978, C2 => 
                           MEM_IN(30), A => n7104, ZN => n7103);
   U7729 : OAI22_X1 port map( A1 => n11375, A2 => n216, B1 => n5171, B2 => n146
                           , ZN => n7104);
   U7730 : AOI22_X1 port map( A1 => n6981, A2 => n5172, B1 => n6982, B2 => 
                           n5173, ZN => n7102);
   U7731 : AOI22_X1 port map( A1 => n6983, A2 => n5174, B1 => n6984, B2 => 
                           n5175, ZN => n7101);
   U7732 : NAND3_X1 port map( A1 => n7105, A2 => n7106, A3 => n7107, ZN => 
                           n12737);
   U7733 : AOI221_X1 port map( B1 => n6977, B2 => n5179, C1 => n6978, C2 => 
                           MEM_IN(31), A => n7108, ZN => n7107);
   U7734 : OAI22_X1 port map( A1 => n11374, A2 => n216, B1 => n5181, B2 => n146
                           , ZN => n7108);
   U7735 : AOI22_X1 port map( A1 => n6981, A2 => n5191, B1 => n6982, B2 => 
                           n5192, ZN => n7106);
   U7736 : AOI22_X1 port map( A1 => n6983, A2 => n5195, B1 => n6984, B2 => 
                           n5196, ZN => n7105);
   U7737 : OAI22_X1 port map( A1 => n7110, A2 => n7114, B1 => n208, B2 => n215,
                           ZN => n7112);
   U7738 : INV_X1 port map( A => n7109, ZN => n7114);
   U7739 : NOR3_X1 port map( A1 => n4841, A2 => n215, A3 => n6077, ZN => n7109)
                           ;
   U7740 : OAI22_X1 port map( A1 => n4786, A2 => n7115, B1 => n7116, B2 => 
                           n5204, ZN => n6980);
   U7741 : NOR2_X1 port map( A1 => n6077, A2 => n7110, ZN => n7116);
   U7742 : NAND2_X1 port map( A1 => n7117, A2 => n6676, ZN => n6077);
   U7743 : INV_X1 port map( A => n6968, ZN => n6676);
   U7744 : INV_X1 port map( A => n7118, ZN => n7115);
   U7745 : OAI211_X1 port map( C1 => n6971, C2 => n5923, A => n7111, B => n5368
                           , ZN => n7118);
   U7746 : AOI21_X1 port map( B1 => n6968, B2 => n5206, A => n7113, ZN => n7111
                           );
   U7747 : NAND2_X1 port map( A1 => n6526, A2 => n6530, ZN => n6968);
   U7748 : AND2_X1 port map( A1 => n6380, A2 => n6227, ZN => n6526);
   U7749 : NAND2_X1 port map( A1 => n7119, A2 => n7120, ZN => n7110);
   U7750 : NOR2_X1 port map( A1 => n6227, A2 => n4787, ZN => n6672);
   U7751 : NAND2_X1 port map( A1 => n5926, A2 => n6531, ZN => n6227);
   U7752 : NAND3_X1 port map( A1 => n7121, A2 => n7122, A3 => n7123, ZN => 
                           n12736);
   U7753 : AOI221_X1 port map( B1 => n7124, B2 => n4863, C1 => n191, C2 => 
                           MEM_IN(0), A => n7125, ZN => n7123);
   U7754 : OAI22_X1 port map( A1 => n11373, A2 => n295, B1 => n4867, B2 => n147
                           , ZN => n7125);
   U7755 : AOI22_X1 port map( A1 => n7127, A2 => n4869, B1 => n7128, B2 => 
                           n4871, ZN => n7122);
   U7756 : AOI22_X1 port map( A1 => n7129, A2 => n4873, B1 => n7130, B2 => 
                           n4875, ZN => n7121);
   U7757 : NAND3_X1 port map( A1 => n7131, A2 => n7132, A3 => n7133, ZN => 
                           n12735);
   U7758 : AOI221_X1 port map( B1 => n7124, B2 => n4879, C1 => n191, C2 => 
                           MEM_IN(1), A => n7134, ZN => n7133);
   U7759 : OAI22_X1 port map( A1 => n11372, A2 => n295, B1 => n4881, B2 => n147
                           , ZN => n7134);
   U7760 : AOI22_X1 port map( A1 => n7127, A2 => n4882, B1 => n7128, B2 => 
                           n4883, ZN => n7132);
   U7761 : AOI22_X1 port map( A1 => n7129, A2 => n4884, B1 => n7130, B2 => 
                           n4885, ZN => n7131);
   U7762 : NAND3_X1 port map( A1 => n7135, A2 => n7136, A3 => n7137, ZN => 
                           n12734);
   U7763 : AOI221_X1 port map( B1 => n7124, B2 => n4889, C1 => n191, C2 => 
                           MEM_IN(2), A => n7138, ZN => n7137);
   U7764 : OAI22_X1 port map( A1 => n11371, A2 => n295, B1 => n4891, B2 => n147
                           , ZN => n7138);
   U7765 : AOI22_X1 port map( A1 => n7127, A2 => n4892, B1 => n7128, B2 => 
                           n4893, ZN => n7136);
   U7766 : AOI22_X1 port map( A1 => n7129, A2 => n4894, B1 => n7130, B2 => 
                           n4895, ZN => n7135);
   U7767 : NAND3_X1 port map( A1 => n7139, A2 => n7140, A3 => n7141, ZN => 
                           n12733);
   U7768 : AOI221_X1 port map( B1 => n7124, B2 => n4899, C1 => n191, C2 => 
                           MEM_IN(3), A => n7142, ZN => n7141);
   U7769 : OAI22_X1 port map( A1 => n11370, A2 => n295, B1 => n4901, B2 => n147
                           , ZN => n7142);
   U7770 : AOI22_X1 port map( A1 => n7127, A2 => n4902, B1 => n7128, B2 => 
                           n4903, ZN => n7140);
   U7771 : AOI22_X1 port map( A1 => n7129, A2 => n4904, B1 => n7130, B2 => 
                           n4905, ZN => n7139);
   U7772 : NAND3_X1 port map( A1 => n7143, A2 => n7144, A3 => n7145, ZN => 
                           n12732);
   U7773 : AOI221_X1 port map( B1 => n7124, B2 => n4909, C1 => n191, C2 => 
                           MEM_IN(4), A => n7146, ZN => n7145);
   U7774 : OAI22_X1 port map( A1 => n11369, A2 => n295, B1 => n4911, B2 => n147
                           , ZN => n7146);
   U7775 : AOI22_X1 port map( A1 => n7127, A2 => n4912, B1 => n7128, B2 => 
                           n4913, ZN => n7144);
   U7776 : AOI22_X1 port map( A1 => n7129, A2 => n4914, B1 => n7130, B2 => 
                           n4915, ZN => n7143);
   U7777 : NAND3_X1 port map( A1 => n7147, A2 => n7148, A3 => n7149, ZN => 
                           n12731);
   U7778 : AOI221_X1 port map( B1 => n7124, B2 => n4919, C1 => n191, C2 => 
                           MEM_IN(5), A => n7150, ZN => n7149);
   U7779 : OAI22_X1 port map( A1 => n11368, A2 => n295, B1 => n4921, B2 => n147
                           , ZN => n7150);
   U7780 : AOI22_X1 port map( A1 => n7127, A2 => n4922, B1 => n7128, B2 => 
                           n4923, ZN => n7148);
   U7781 : AOI22_X1 port map( A1 => n7129, A2 => n4924, B1 => n7130, B2 => 
                           n4925, ZN => n7147);
   U7782 : NAND3_X1 port map( A1 => n7151, A2 => n7152, A3 => n7153, ZN => 
                           n12730);
   U7783 : AOI221_X1 port map( B1 => n7124, B2 => n4929, C1 => n191, C2 => 
                           MEM_IN(6), A => n7154, ZN => n7153);
   U7784 : OAI22_X1 port map( A1 => n11367, A2 => n295, B1 => n4931, B2 => n147
                           , ZN => n7154);
   U7785 : AOI22_X1 port map( A1 => n7127, A2 => n4932, B1 => n7128, B2 => 
                           n4933, ZN => n7152);
   U7786 : AOI22_X1 port map( A1 => n7129, A2 => n4934, B1 => n7130, B2 => 
                           n4935, ZN => n7151);
   U7787 : NAND3_X1 port map( A1 => n7155, A2 => n7156, A3 => n7157, ZN => 
                           n12729);
   U7788 : AOI221_X1 port map( B1 => n7124, B2 => n4939, C1 => n191, C2 => 
                           MEM_IN(7), A => n7158, ZN => n7157);
   U7789 : OAI22_X1 port map( A1 => n11366, A2 => n295, B1 => n4941, B2 => n147
                           , ZN => n7158);
   U7790 : AOI22_X1 port map( A1 => n7127, A2 => n4942, B1 => n7128, B2 => 
                           n4943, ZN => n7156);
   U7791 : AOI22_X1 port map( A1 => n7129, A2 => n4944, B1 => n7130, B2 => 
                           n4945, ZN => n7155);
   U7792 : NAND3_X1 port map( A1 => n7159, A2 => n7160, A3 => n7161, ZN => 
                           n12728);
   U7793 : AOI221_X1 port map( B1 => n7124, B2 => n4949, C1 => n191, C2 => 
                           MEM_IN(8), A => n7162, ZN => n7161);
   U7794 : OAI22_X1 port map( A1 => n11365, A2 => n295, B1 => n4951, B2 => n147
                           , ZN => n7162);
   U7795 : AOI22_X1 port map( A1 => n7127, A2 => n4952, B1 => n7128, B2 => 
                           n4953, ZN => n7160);
   U7796 : AOI22_X1 port map( A1 => n7129, A2 => n4954, B1 => n7130, B2 => 
                           n4955, ZN => n7159);
   U7797 : NAND3_X1 port map( A1 => n7163, A2 => n7164, A3 => n7165, ZN => 
                           n12727);
   U7798 : AOI221_X1 port map( B1 => n7124, B2 => n4959, C1 => n191, C2 => 
                           MEM_IN(9), A => n7166, ZN => n7165);
   U7799 : OAI22_X1 port map( A1 => n11364, A2 => n295, B1 => n4961, B2 => n147
                           , ZN => n7166);
   U7800 : AOI22_X1 port map( A1 => n7127, A2 => n4962, B1 => n7128, B2 => 
                           n4963, ZN => n7164);
   U7801 : AOI22_X1 port map( A1 => n7129, A2 => n4964, B1 => n7130, B2 => 
                           n4965, ZN => n7163);
   U7802 : NAND3_X1 port map( A1 => n7167, A2 => n7168, A3 => n7169, ZN => 
                           n12726);
   U7803 : AOI221_X1 port map( B1 => n7124, B2 => n4969, C1 => n191, C2 => 
                           MEM_IN(10), A => n7170, ZN => n7169);
   U7804 : OAI22_X1 port map( A1 => n11363, A2 => n295, B1 => n4971, B2 => n147
                           , ZN => n7170);
   U7805 : AOI22_X1 port map( A1 => n7127, A2 => n4972, B1 => n7128, B2 => 
                           n4973, ZN => n7168);
   U7806 : AOI22_X1 port map( A1 => n7129, A2 => n4974, B1 => n7130, B2 => 
                           n4975, ZN => n7167);
   U7807 : NAND3_X1 port map( A1 => n7171, A2 => n7172, A3 => n7173, ZN => 
                           n12725);
   U7808 : AOI221_X1 port map( B1 => n7124, B2 => n4979, C1 => n191, C2 => 
                           MEM_IN(11), A => n7174, ZN => n7173);
   U7809 : OAI22_X1 port map( A1 => n11362, A2 => n295, B1 => n4981, B2 => n147
                           , ZN => n7174);
   U7810 : AOI22_X1 port map( A1 => n7127, A2 => n4982, B1 => n7128, B2 => 
                           n4983, ZN => n7172);
   U7811 : AOI22_X1 port map( A1 => n7129, A2 => n4984, B1 => n7130, B2 => 
                           n4985, ZN => n7171);
   U7812 : NAND3_X1 port map( A1 => n7175, A2 => n7176, A3 => n7177, ZN => 
                           n12724);
   U7813 : AOI221_X1 port map( B1 => n7124, B2 => n4989, C1 => n191, C2 => 
                           MEM_IN(12), A => n7178, ZN => n7177);
   U7814 : OAI22_X1 port map( A1 => n11361, A2 => n295, B1 => n4991, B2 => n147
                           , ZN => n7178);
   U7815 : AOI22_X1 port map( A1 => n7127, A2 => n4992, B1 => n7128, B2 => 
                           n4993, ZN => n7176);
   U7816 : AOI22_X1 port map( A1 => n7129, A2 => n4994, B1 => n7130, B2 => 
                           n4995, ZN => n7175);
   U7817 : NAND3_X1 port map( A1 => n7179, A2 => n7180, A3 => n7181, ZN => 
                           n12723);
   U7818 : AOI221_X1 port map( B1 => n7124, B2 => n4999, C1 => n191, C2 => 
                           MEM_IN(13), A => n7182, ZN => n7181);
   U7819 : OAI22_X1 port map( A1 => n11360, A2 => n295, B1 => n5001, B2 => n147
                           , ZN => n7182);
   U7820 : AOI22_X1 port map( A1 => n7127, A2 => n5002, B1 => n7128, B2 => 
                           n5003, ZN => n7180);
   U7821 : AOI22_X1 port map( A1 => n7129, A2 => n5004, B1 => n7130, B2 => 
                           n5005, ZN => n7179);
   U7822 : NAND3_X1 port map( A1 => n7183, A2 => n7184, A3 => n7185, ZN => 
                           n12722);
   U7823 : AOI221_X1 port map( B1 => n7124, B2 => n5009, C1 => n191, C2 => 
                           MEM_IN(14), A => n7186, ZN => n7185);
   U7824 : OAI22_X1 port map( A1 => n11359, A2 => n295, B1 => n5011, B2 => n147
                           , ZN => n7186);
   U7825 : AOI22_X1 port map( A1 => n7127, A2 => n5012, B1 => n7128, B2 => 
                           n5013, ZN => n7184);
   U7826 : AOI22_X1 port map( A1 => n7129, A2 => n5014, B1 => n7130, B2 => 
                           n5015, ZN => n7183);
   U7827 : NAND3_X1 port map( A1 => n7187, A2 => n7188, A3 => n7189, ZN => 
                           n12721);
   U7828 : AOI221_X1 port map( B1 => n7124, B2 => n5019, C1 => n191, C2 => 
                           MEM_IN(15), A => n7190, ZN => n7189);
   U7829 : OAI22_X1 port map( A1 => n11358, A2 => n295, B1 => n5021, B2 => n147
                           , ZN => n7190);
   U7830 : AOI22_X1 port map( A1 => n7127, A2 => n5022, B1 => n7128, B2 => 
                           n5023, ZN => n7188);
   U7831 : AOI22_X1 port map( A1 => n7129, A2 => n5024, B1 => n7130, B2 => 
                           n5025, ZN => n7187);
   U7832 : NAND3_X1 port map( A1 => n7191, A2 => n7192, A3 => n7193, ZN => 
                           n12720);
   U7833 : AOI221_X1 port map( B1 => n7124, B2 => n5029, C1 => n191, C2 => 
                           MEM_IN(16), A => n7194, ZN => n7193);
   U7834 : OAI22_X1 port map( A1 => n11357, A2 => n295, B1 => n5031, B2 => n147
                           , ZN => n7194);
   U7835 : AOI22_X1 port map( A1 => n7127, A2 => n5032, B1 => n7128, B2 => 
                           n5033, ZN => n7192);
   U7836 : AOI22_X1 port map( A1 => n7129, A2 => n5034, B1 => n7130, B2 => 
                           n5035, ZN => n7191);
   U7837 : NAND3_X1 port map( A1 => n7195, A2 => n7196, A3 => n7197, ZN => 
                           n12719);
   U7838 : AOI221_X1 port map( B1 => n7124, B2 => n5039, C1 => n191, C2 => 
                           MEM_IN(17), A => n7198, ZN => n7197);
   U7839 : OAI22_X1 port map( A1 => n11356, A2 => n295, B1 => n5041, B2 => n147
                           , ZN => n7198);
   U7840 : AOI22_X1 port map( A1 => n7127, A2 => n5042, B1 => n7128, B2 => 
                           n5043, ZN => n7196);
   U7841 : AOI22_X1 port map( A1 => n7129, A2 => n5044, B1 => n7130, B2 => 
                           n5045, ZN => n7195);
   U7842 : NAND3_X1 port map( A1 => n7199, A2 => n7200, A3 => n7201, ZN => 
                           n12718);
   U7843 : AOI221_X1 port map( B1 => n7124, B2 => n5049, C1 => n191, C2 => 
                           MEM_IN(18), A => n7202, ZN => n7201);
   U7844 : OAI22_X1 port map( A1 => n11355, A2 => n295, B1 => n5051, B2 => n147
                           , ZN => n7202);
   U7845 : AOI22_X1 port map( A1 => n7127, A2 => n5052, B1 => n7128, B2 => 
                           n5053, ZN => n7200);
   U7846 : AOI22_X1 port map( A1 => n7129, A2 => n5054, B1 => n7130, B2 => 
                           n5055, ZN => n7199);
   U7847 : NAND3_X1 port map( A1 => n7203, A2 => n7204, A3 => n7205, ZN => 
                           n12717);
   U7848 : AOI221_X1 port map( B1 => n7124, B2 => n5059, C1 => n191, C2 => 
                           MEM_IN(19), A => n7206, ZN => n7205);
   U7849 : OAI22_X1 port map( A1 => n11354, A2 => n295, B1 => n5061, B2 => n147
                           , ZN => n7206);
   U7850 : AOI22_X1 port map( A1 => n7127, A2 => n5062, B1 => n7128, B2 => 
                           n5063, ZN => n7204);
   U7851 : AOI22_X1 port map( A1 => n7129, A2 => n5064, B1 => n7130, B2 => 
                           n5065, ZN => n7203);
   U7852 : NAND3_X1 port map( A1 => n7207, A2 => n7208, A3 => n7209, ZN => 
                           n12716);
   U7853 : AOI221_X1 port map( B1 => n7124, B2 => n5069, C1 => n191, C2 => 
                           MEM_IN(20), A => n7210, ZN => n7209);
   U7854 : OAI22_X1 port map( A1 => n11353, A2 => n295, B1 => n5071, B2 => n147
                           , ZN => n7210);
   U7855 : AOI22_X1 port map( A1 => n7127, A2 => n5072, B1 => n7128, B2 => 
                           n5073, ZN => n7208);
   U7856 : AOI22_X1 port map( A1 => n7129, A2 => n5074, B1 => n7130, B2 => 
                           n5075, ZN => n7207);
   U7857 : NAND3_X1 port map( A1 => n7211, A2 => n7212, A3 => n7213, ZN => 
                           n12715);
   U7858 : AOI221_X1 port map( B1 => n7124, B2 => n5079, C1 => n191, C2 => 
                           MEM_IN(21), A => n7214, ZN => n7213);
   U7859 : OAI22_X1 port map( A1 => n11352, A2 => n295, B1 => n5081, B2 => n147
                           , ZN => n7214);
   U7860 : AOI22_X1 port map( A1 => n7127, A2 => n5082, B1 => n7128, B2 => 
                           n5083, ZN => n7212);
   U7861 : AOI22_X1 port map( A1 => n7129, A2 => n5084, B1 => n7130, B2 => 
                           n5085, ZN => n7211);
   U7862 : NAND3_X1 port map( A1 => n7215, A2 => n7216, A3 => n7217, ZN => 
                           n12714);
   U7863 : AOI221_X1 port map( B1 => n7124, B2 => n5089, C1 => n191, C2 => 
                           MEM_IN(22), A => n7218, ZN => n7217);
   U7864 : OAI22_X1 port map( A1 => n11351, A2 => n295, B1 => n5091, B2 => n147
                           , ZN => n7218);
   U7865 : AOI22_X1 port map( A1 => n7127, A2 => n5092, B1 => n7128, B2 => 
                           n5093, ZN => n7216);
   U7866 : AOI22_X1 port map( A1 => n7129, A2 => n5094, B1 => n7130, B2 => 
                           n5095, ZN => n7215);
   U7867 : NAND3_X1 port map( A1 => n7219, A2 => n7220, A3 => n7221, ZN => 
                           n12713);
   U7868 : AOI221_X1 port map( B1 => n7124, B2 => n5099, C1 => n191, C2 => 
                           MEM_IN(23), A => n7222, ZN => n7221);
   U7869 : OAI22_X1 port map( A1 => n11350, A2 => n295, B1 => n5101, B2 => n147
                           , ZN => n7222);
   U7870 : AOI22_X1 port map( A1 => n7127, A2 => n5102, B1 => n7128, B2 => 
                           n5103, ZN => n7220);
   U7871 : AOI22_X1 port map( A1 => n7129, A2 => n5104, B1 => n7130, B2 => 
                           n5105, ZN => n7219);
   U7872 : NAND3_X1 port map( A1 => n7223, A2 => n7224, A3 => n7225, ZN => 
                           n12712);
   U7873 : AOI221_X1 port map( B1 => n7124, B2 => n5109, C1 => n191, C2 => 
                           MEM_IN(24), A => n7226, ZN => n7225);
   U7874 : OAI22_X1 port map( A1 => n11349, A2 => n295, B1 => n5111, B2 => n147
                           , ZN => n7226);
   U7875 : AOI22_X1 port map( A1 => n7127, A2 => n5112, B1 => n7128, B2 => 
                           n5113, ZN => n7224);
   U7876 : AOI22_X1 port map( A1 => n7129, A2 => n5114, B1 => n7130, B2 => 
                           n5115, ZN => n7223);
   U7877 : NAND3_X1 port map( A1 => n7227, A2 => n7228, A3 => n7229, ZN => 
                           n12711);
   U7878 : AOI221_X1 port map( B1 => n7124, B2 => n5119, C1 => n191, C2 => 
                           MEM_IN(25), A => n7230, ZN => n7229);
   U7879 : OAI22_X1 port map( A1 => n11348, A2 => n295, B1 => n5121, B2 => n147
                           , ZN => n7230);
   U7880 : AOI22_X1 port map( A1 => n7127, A2 => n5122, B1 => n7128, B2 => 
                           n5123, ZN => n7228);
   U7881 : AOI22_X1 port map( A1 => n7129, A2 => n5124, B1 => n7130, B2 => 
                           n5125, ZN => n7227);
   U7882 : NAND3_X1 port map( A1 => n7231, A2 => n7232, A3 => n7233, ZN => 
                           n12710);
   U7883 : AOI221_X1 port map( B1 => n7124, B2 => n5129, C1 => n191, C2 => 
                           MEM_IN(26), A => n7234, ZN => n7233);
   U7884 : OAI22_X1 port map( A1 => n11347, A2 => n295, B1 => n5131, B2 => n147
                           , ZN => n7234);
   U7885 : AOI22_X1 port map( A1 => n7127, A2 => n5132, B1 => n7128, B2 => 
                           n5133, ZN => n7232);
   U7886 : AOI22_X1 port map( A1 => n7129, A2 => n5134, B1 => n7130, B2 => 
                           n5135, ZN => n7231);
   U7887 : NAND3_X1 port map( A1 => n7235, A2 => n7236, A3 => n7237, ZN => 
                           n12709);
   U7888 : AOI221_X1 port map( B1 => n7124, B2 => n5139, C1 => n191, C2 => 
                           MEM_IN(27), A => n7238, ZN => n7237);
   U7889 : OAI22_X1 port map( A1 => n11346, A2 => n295, B1 => n5141, B2 => n147
                           , ZN => n7238);
   U7890 : AOI22_X1 port map( A1 => n7127, A2 => n5142, B1 => n7128, B2 => 
                           n5143, ZN => n7236);
   U7891 : AOI22_X1 port map( A1 => n7129, A2 => n5144, B1 => n7130, B2 => 
                           n5145, ZN => n7235);
   U7892 : NAND3_X1 port map( A1 => n7239, A2 => n7240, A3 => n7241, ZN => 
                           n12708);
   U7893 : AOI221_X1 port map( B1 => n7124, B2 => n5149, C1 => n191, C2 => 
                           MEM_IN(28), A => n7242, ZN => n7241);
   U7894 : OAI22_X1 port map( A1 => n11345, A2 => n295, B1 => n5151, B2 => n147
                           , ZN => n7242);
   U7895 : AOI22_X1 port map( A1 => n7127, A2 => n5152, B1 => n7128, B2 => 
                           n5153, ZN => n7240);
   U7896 : AOI22_X1 port map( A1 => n7129, A2 => n5154, B1 => n7130, B2 => 
                           n5155, ZN => n7239);
   U7897 : NAND3_X1 port map( A1 => n7243, A2 => n7244, A3 => n7245, ZN => 
                           n12707);
   U7898 : AOI221_X1 port map( B1 => n7124, B2 => n5159, C1 => n191, C2 => 
                           MEM_IN(29), A => n7246, ZN => n7245);
   U7899 : OAI22_X1 port map( A1 => n11344, A2 => n295, B1 => n5161, B2 => n147
                           , ZN => n7246);
   U7900 : AOI22_X1 port map( A1 => n7127, A2 => n5162, B1 => n7128, B2 => 
                           n5163, ZN => n7244);
   U7901 : AOI22_X1 port map( A1 => n7129, A2 => n5164, B1 => n7130, B2 => 
                           n5165, ZN => n7243);
   U7902 : NAND3_X1 port map( A1 => n7247, A2 => n7248, A3 => n7249, ZN => 
                           n12706);
   U7903 : AOI221_X1 port map( B1 => n7124, B2 => n5169, C1 => n191, C2 => 
                           MEM_IN(30), A => n7250, ZN => n7249);
   U7904 : OAI22_X1 port map( A1 => n11343, A2 => n295, B1 => n5171, B2 => n147
                           , ZN => n7250);
   U7905 : AOI22_X1 port map( A1 => n7127, A2 => n5172, B1 => n7128, B2 => 
                           n5173, ZN => n7248);
   U7906 : AOI22_X1 port map( A1 => n7129, A2 => n5174, B1 => n7130, B2 => 
                           n5175, ZN => n7247);
   U7907 : NAND3_X1 port map( A1 => n7251, A2 => n7252, A3 => n7253, ZN => 
                           n12705);
   U7908 : AOI221_X1 port map( B1 => n7124, B2 => n5179, C1 => n191, C2 => 
                           MEM_IN(31), A => n7254, ZN => n7253);
   U7909 : OAI22_X1 port map( A1 => n11342, A2 => n295, B1 => n5181, B2 => n147
                           , ZN => n7254);
   U7910 : INV_X1 port map( A => n7258, ZN => n7257);
   U7911 : AOI22_X1 port map( A1 => n7127, A2 => n5191, B1 => n7128, B2 => 
                           n5192, ZN => n7252);
   U7912 : AOI22_X1 port map( A1 => n7129, A2 => n5195, B1 => n7130, B2 => 
                           n5196, ZN => n7251);
   U7913 : OAI22_X1 port map( A1 => n7258, A2 => n7256, B1 => n208, B2 => n294,
                           ZN => n7259);
   U7914 : NAND3_X1 port map( A1 => n208, A2 => n295, A3 => n6226, ZN => n7256)
                           ;
   U7915 : INV_X1 port map( A => n7255, ZN => n6226);
   U7916 : OAI22_X1 port map( A1 => n4786, A2 => n7262, B1 => n7263, B2 => 
                           n5204, ZN => n7126);
   U7917 : NOR2_X1 port map( A1 => n7255, A2 => n7258, ZN => n7263);
   U7918 : NAND4_X1 port map( A1 => n7117, A2 => n7120, A3 => n6530, A4 => 
                           n6380, ZN => n7255);
   U7919 : NOR4_X1 port map( A1 => n7264, A2 => n7113, A3 => RESET, A4 => n7261
                           , ZN => n7262);
   U7920 : OAI211_X1 port map( C1 => n6076, C2 => n6971, A => n6815, B => n6961
                           , ZN => n7264);
   U7921 : INV_X1 port map( A => n6963, ZN => n6815);
   U7922 : NAND2_X1 port map( A1 => n7265, A2 => n7266, ZN => n7258);
   U7923 : NOR2_X1 port map( A1 => n6380, A2 => n4787, ZN => n6963);
   U7924 : NAND2_X1 port map( A1 => n6079, A2 => n6531, ZN => n6380);
   U7925 : NAND3_X1 port map( A1 => n7267, A2 => n7268, A3 => n7269, ZN => 
                           n12704);
   U7926 : AOI221_X1 port map( B1 => n7270, B2 => n4863, C1 => n192, C2 => 
                           MEM_IN(0), A => n7271, ZN => n7269);
   U7927 : OAI22_X1 port map( A1 => n11341, A2 => n297, B1 => n4867, B2 => n144
                           , ZN => n7271);
   U7928 : AOI22_X1 port map( A1 => n7273, A2 => n4869, B1 => n7274, B2 => 
                           n4871, ZN => n7268);
   U7929 : AOI22_X1 port map( A1 => n7275, A2 => n4873, B1 => n7276, B2 => 
                           n4875, ZN => n7267);
   U7930 : NAND3_X1 port map( A1 => n7277, A2 => n7278, A3 => n7279, ZN => 
                           n12703);
   U7931 : AOI221_X1 port map( B1 => n7270, B2 => n4879, C1 => n192, C2 => 
                           MEM_IN(1), A => n7280, ZN => n7279);
   U7932 : OAI22_X1 port map( A1 => n11340, A2 => n297, B1 => n4881, B2 => n144
                           , ZN => n7280);
   U7933 : AOI22_X1 port map( A1 => n7273, A2 => n4882, B1 => n7274, B2 => 
                           n4883, ZN => n7278);
   U7934 : AOI22_X1 port map( A1 => n7275, A2 => n4884, B1 => n7276, B2 => 
                           n4885, ZN => n7277);
   U7935 : NAND3_X1 port map( A1 => n7281, A2 => n7282, A3 => n7283, ZN => 
                           n12702);
   U7936 : AOI221_X1 port map( B1 => n7270, B2 => n4889, C1 => n192, C2 => 
                           MEM_IN(2), A => n7284, ZN => n7283);
   U7937 : OAI22_X1 port map( A1 => n11339, A2 => n297, B1 => n4891, B2 => n144
                           , ZN => n7284);
   U7938 : AOI22_X1 port map( A1 => n7273, A2 => n4892, B1 => n7274, B2 => 
                           n4893, ZN => n7282);
   U7939 : AOI22_X1 port map( A1 => n7275, A2 => n4894, B1 => n7276, B2 => 
                           n4895, ZN => n7281);
   U7940 : NAND3_X1 port map( A1 => n7285, A2 => n7286, A3 => n7287, ZN => 
                           n12701);
   U7941 : AOI221_X1 port map( B1 => n7270, B2 => n4899, C1 => n192, C2 => 
                           MEM_IN(3), A => n7288, ZN => n7287);
   U7942 : OAI22_X1 port map( A1 => n11338, A2 => n297, B1 => n4901, B2 => n144
                           , ZN => n7288);
   U7943 : AOI22_X1 port map( A1 => n7273, A2 => n4902, B1 => n7274, B2 => 
                           n4903, ZN => n7286);
   U7944 : AOI22_X1 port map( A1 => n7275, A2 => n4904, B1 => n7276, B2 => 
                           n4905, ZN => n7285);
   U7945 : NAND3_X1 port map( A1 => n7289, A2 => n7290, A3 => n7291, ZN => 
                           n12700);
   U7946 : AOI221_X1 port map( B1 => n7270, B2 => n4909, C1 => n192, C2 => 
                           MEM_IN(4), A => n7292, ZN => n7291);
   U7947 : OAI22_X1 port map( A1 => n11337, A2 => n297, B1 => n4911, B2 => n144
                           , ZN => n7292);
   U7948 : AOI22_X1 port map( A1 => n7273, A2 => n4912, B1 => n7274, B2 => 
                           n4913, ZN => n7290);
   U7949 : AOI22_X1 port map( A1 => n7275, A2 => n4914, B1 => n7276, B2 => 
                           n4915, ZN => n7289);
   U7950 : NAND3_X1 port map( A1 => n7293, A2 => n7294, A3 => n7295, ZN => 
                           n12699);
   U7951 : AOI221_X1 port map( B1 => n7270, B2 => n4919, C1 => n192, C2 => 
                           MEM_IN(5), A => n7296, ZN => n7295);
   U7952 : OAI22_X1 port map( A1 => n11336, A2 => n297, B1 => n4921, B2 => n144
                           , ZN => n7296);
   U7953 : AOI22_X1 port map( A1 => n7273, A2 => n4922, B1 => n7274, B2 => 
                           n4923, ZN => n7294);
   U7954 : AOI22_X1 port map( A1 => n7275, A2 => n4924, B1 => n7276, B2 => 
                           n4925, ZN => n7293);
   U7955 : NAND3_X1 port map( A1 => n7297, A2 => n7298, A3 => n7299, ZN => 
                           n12698);
   U7956 : AOI221_X1 port map( B1 => n7270, B2 => n4929, C1 => n192, C2 => 
                           MEM_IN(6), A => n7300, ZN => n7299);
   U7957 : OAI22_X1 port map( A1 => n11335, A2 => n297, B1 => n4931, B2 => n144
                           , ZN => n7300);
   U7958 : AOI22_X1 port map( A1 => n7273, A2 => n4932, B1 => n7274, B2 => 
                           n4933, ZN => n7298);
   U7959 : AOI22_X1 port map( A1 => n7275, A2 => n4934, B1 => n7276, B2 => 
                           n4935, ZN => n7297);
   U7960 : NAND3_X1 port map( A1 => n7301, A2 => n7302, A3 => n7303, ZN => 
                           n12697);
   U7961 : AOI221_X1 port map( B1 => n7270, B2 => n4939, C1 => n192, C2 => 
                           MEM_IN(7), A => n7304, ZN => n7303);
   U7962 : OAI22_X1 port map( A1 => n11334, A2 => n297, B1 => n4941, B2 => n144
                           , ZN => n7304);
   U7963 : AOI22_X1 port map( A1 => n7273, A2 => n4942, B1 => n7274, B2 => 
                           n4943, ZN => n7302);
   U7964 : AOI22_X1 port map( A1 => n7275, A2 => n4944, B1 => n7276, B2 => 
                           n4945, ZN => n7301);
   U7965 : NAND3_X1 port map( A1 => n7305, A2 => n7306, A3 => n7307, ZN => 
                           n12696);
   U7966 : AOI221_X1 port map( B1 => n7270, B2 => n4949, C1 => n192, C2 => 
                           MEM_IN(8), A => n7308, ZN => n7307);
   U7967 : OAI22_X1 port map( A1 => n11333, A2 => n297, B1 => n4951, B2 => n144
                           , ZN => n7308);
   U7968 : AOI22_X1 port map( A1 => n7273, A2 => n4952, B1 => n7274, B2 => 
                           n4953, ZN => n7306);
   U7969 : AOI22_X1 port map( A1 => n7275, A2 => n4954, B1 => n7276, B2 => 
                           n4955, ZN => n7305);
   U7970 : NAND3_X1 port map( A1 => n7309, A2 => n7310, A3 => n7311, ZN => 
                           n12695);
   U7971 : AOI221_X1 port map( B1 => n7270, B2 => n4959, C1 => n192, C2 => 
                           MEM_IN(9), A => n7312, ZN => n7311);
   U7972 : OAI22_X1 port map( A1 => n11332, A2 => n297, B1 => n4961, B2 => n144
                           , ZN => n7312);
   U7973 : AOI22_X1 port map( A1 => n7273, A2 => n4962, B1 => n7274, B2 => 
                           n4963, ZN => n7310);
   U7974 : AOI22_X1 port map( A1 => n7275, A2 => n4964, B1 => n7276, B2 => 
                           n4965, ZN => n7309);
   U7975 : NAND3_X1 port map( A1 => n7313, A2 => n7314, A3 => n7315, ZN => 
                           n12694);
   U7976 : AOI221_X1 port map( B1 => n7270, B2 => n4969, C1 => n192, C2 => 
                           MEM_IN(10), A => n7316, ZN => n7315);
   U7977 : OAI22_X1 port map( A1 => n11331, A2 => n297, B1 => n4971, B2 => n144
                           , ZN => n7316);
   U7978 : AOI22_X1 port map( A1 => n7273, A2 => n4972, B1 => n7274, B2 => 
                           n4973, ZN => n7314);
   U7979 : AOI22_X1 port map( A1 => n7275, A2 => n4974, B1 => n7276, B2 => 
                           n4975, ZN => n7313);
   U7980 : NAND3_X1 port map( A1 => n7317, A2 => n7318, A3 => n7319, ZN => 
                           n12693);
   U7981 : AOI221_X1 port map( B1 => n7270, B2 => n4979, C1 => n192, C2 => 
                           MEM_IN(11), A => n7320, ZN => n7319);
   U7982 : OAI22_X1 port map( A1 => n11330, A2 => n297, B1 => n4981, B2 => n144
                           , ZN => n7320);
   U7983 : AOI22_X1 port map( A1 => n7273, A2 => n4982, B1 => n7274, B2 => 
                           n4983, ZN => n7318);
   U7984 : AOI22_X1 port map( A1 => n7275, A2 => n4984, B1 => n7276, B2 => 
                           n4985, ZN => n7317);
   U7985 : NAND3_X1 port map( A1 => n7321, A2 => n7322, A3 => n7323, ZN => 
                           n12692);
   U7986 : AOI221_X1 port map( B1 => n7270, B2 => n4989, C1 => n192, C2 => 
                           MEM_IN(12), A => n7324, ZN => n7323);
   U7987 : OAI22_X1 port map( A1 => n11329, A2 => n297, B1 => n4991, B2 => n144
                           , ZN => n7324);
   U7988 : AOI22_X1 port map( A1 => n7273, A2 => n4992, B1 => n7274, B2 => 
                           n4993, ZN => n7322);
   U7989 : AOI22_X1 port map( A1 => n7275, A2 => n4994, B1 => n7276, B2 => 
                           n4995, ZN => n7321);
   U7990 : NAND3_X1 port map( A1 => n7325, A2 => n7326, A3 => n7327, ZN => 
                           n12691);
   U7991 : AOI221_X1 port map( B1 => n7270, B2 => n4999, C1 => n192, C2 => 
                           MEM_IN(13), A => n7328, ZN => n7327);
   U7992 : OAI22_X1 port map( A1 => n11328, A2 => n297, B1 => n5001, B2 => n144
                           , ZN => n7328);
   U7993 : AOI22_X1 port map( A1 => n7273, A2 => n5002, B1 => n7274, B2 => 
                           n5003, ZN => n7326);
   U7994 : AOI22_X1 port map( A1 => n7275, A2 => n5004, B1 => n7276, B2 => 
                           n5005, ZN => n7325);
   U7995 : NAND3_X1 port map( A1 => n7329, A2 => n7330, A3 => n7331, ZN => 
                           n12690);
   U7996 : AOI221_X1 port map( B1 => n7270, B2 => n5009, C1 => n192, C2 => 
                           MEM_IN(14), A => n7332, ZN => n7331);
   U7997 : OAI22_X1 port map( A1 => n11327, A2 => n297, B1 => n5011, B2 => n144
                           , ZN => n7332);
   U7998 : AOI22_X1 port map( A1 => n7273, A2 => n5012, B1 => n7274, B2 => 
                           n5013, ZN => n7330);
   U7999 : AOI22_X1 port map( A1 => n7275, A2 => n5014, B1 => n7276, B2 => 
                           n5015, ZN => n7329);
   U8000 : NAND3_X1 port map( A1 => n7333, A2 => n7334, A3 => n7335, ZN => 
                           n12689);
   U8001 : AOI221_X1 port map( B1 => n7270, B2 => n5019, C1 => n192, C2 => 
                           MEM_IN(15), A => n7336, ZN => n7335);
   U8002 : OAI22_X1 port map( A1 => n11326, A2 => n297, B1 => n5021, B2 => n144
                           , ZN => n7336);
   U8003 : AOI22_X1 port map( A1 => n7273, A2 => n5022, B1 => n7274, B2 => 
                           n5023, ZN => n7334);
   U8004 : AOI22_X1 port map( A1 => n7275, A2 => n5024, B1 => n7276, B2 => 
                           n5025, ZN => n7333);
   U8005 : NAND3_X1 port map( A1 => n7337, A2 => n7338, A3 => n7339, ZN => 
                           n12688);
   U8006 : AOI221_X1 port map( B1 => n7270, B2 => n5029, C1 => n192, C2 => 
                           MEM_IN(16), A => n7340, ZN => n7339);
   U8007 : OAI22_X1 port map( A1 => n11325, A2 => n297, B1 => n5031, B2 => n144
                           , ZN => n7340);
   U8008 : AOI22_X1 port map( A1 => n7273, A2 => n5032, B1 => n7274, B2 => 
                           n5033, ZN => n7338);
   U8009 : AOI22_X1 port map( A1 => n7275, A2 => n5034, B1 => n7276, B2 => 
                           n5035, ZN => n7337);
   U8010 : NAND3_X1 port map( A1 => n7341, A2 => n7342, A3 => n7343, ZN => 
                           n12687);
   U8011 : AOI221_X1 port map( B1 => n7270, B2 => n5039, C1 => n192, C2 => 
                           MEM_IN(17), A => n7344, ZN => n7343);
   U8012 : OAI22_X1 port map( A1 => n11324, A2 => n297, B1 => n5041, B2 => n144
                           , ZN => n7344);
   U8013 : AOI22_X1 port map( A1 => n7273, A2 => n5042, B1 => n7274, B2 => 
                           n5043, ZN => n7342);
   U8014 : AOI22_X1 port map( A1 => n7275, A2 => n5044, B1 => n7276, B2 => 
                           n5045, ZN => n7341);
   U8015 : NAND3_X1 port map( A1 => n7345, A2 => n7346, A3 => n7347, ZN => 
                           n12686);
   U8016 : AOI221_X1 port map( B1 => n7270, B2 => n5049, C1 => n192, C2 => 
                           MEM_IN(18), A => n7348, ZN => n7347);
   U8017 : OAI22_X1 port map( A1 => n11323, A2 => n297, B1 => n5051, B2 => n144
                           , ZN => n7348);
   U8018 : AOI22_X1 port map( A1 => n7273, A2 => n5052, B1 => n7274, B2 => 
                           n5053, ZN => n7346);
   U8019 : AOI22_X1 port map( A1 => n7275, A2 => n5054, B1 => n7276, B2 => 
                           n5055, ZN => n7345);
   U8020 : NAND3_X1 port map( A1 => n7349, A2 => n7350, A3 => n7351, ZN => 
                           n12685);
   U8021 : AOI221_X1 port map( B1 => n7270, B2 => n5059, C1 => n192, C2 => 
                           MEM_IN(19), A => n7352, ZN => n7351);
   U8022 : OAI22_X1 port map( A1 => n11322, A2 => n297, B1 => n5061, B2 => n144
                           , ZN => n7352);
   U8023 : AOI22_X1 port map( A1 => n7273, A2 => n5062, B1 => n7274, B2 => 
                           n5063, ZN => n7350);
   U8024 : AOI22_X1 port map( A1 => n7275, A2 => n5064, B1 => n7276, B2 => 
                           n5065, ZN => n7349);
   U8025 : NAND3_X1 port map( A1 => n7353, A2 => n7354, A3 => n7355, ZN => 
                           n12684);
   U8026 : AOI221_X1 port map( B1 => n7270, B2 => n5069, C1 => n192, C2 => 
                           MEM_IN(20), A => n7356, ZN => n7355);
   U8027 : OAI22_X1 port map( A1 => n11321, A2 => n297, B1 => n5071, B2 => n144
                           , ZN => n7356);
   U8028 : AOI22_X1 port map( A1 => n7273, A2 => n5072, B1 => n7274, B2 => 
                           n5073, ZN => n7354);
   U8029 : AOI22_X1 port map( A1 => n7275, A2 => n5074, B1 => n7276, B2 => 
                           n5075, ZN => n7353);
   U8030 : NAND3_X1 port map( A1 => n7357, A2 => n7358, A3 => n7359, ZN => 
                           n12683);
   U8031 : AOI221_X1 port map( B1 => n7270, B2 => n5079, C1 => n192, C2 => 
                           MEM_IN(21), A => n7360, ZN => n7359);
   U8032 : OAI22_X1 port map( A1 => n11320, A2 => n297, B1 => n5081, B2 => n144
                           , ZN => n7360);
   U8033 : AOI22_X1 port map( A1 => n7273, A2 => n5082, B1 => n7274, B2 => 
                           n5083, ZN => n7358);
   U8034 : AOI22_X1 port map( A1 => n7275, A2 => n5084, B1 => n7276, B2 => 
                           n5085, ZN => n7357);
   U8035 : NAND3_X1 port map( A1 => n7361, A2 => n7362, A3 => n7363, ZN => 
                           n12682);
   U8036 : AOI221_X1 port map( B1 => n7270, B2 => n5089, C1 => n192, C2 => 
                           MEM_IN(22), A => n7364, ZN => n7363);
   U8037 : OAI22_X1 port map( A1 => n11319, A2 => n297, B1 => n5091, B2 => n144
                           , ZN => n7364);
   U8038 : AOI22_X1 port map( A1 => n7273, A2 => n5092, B1 => n7274, B2 => 
                           n5093, ZN => n7362);
   U8039 : AOI22_X1 port map( A1 => n7275, A2 => n5094, B1 => n7276, B2 => 
                           n5095, ZN => n7361);
   U8040 : NAND3_X1 port map( A1 => n7365, A2 => n7366, A3 => n7367, ZN => 
                           n12681);
   U8041 : AOI221_X1 port map( B1 => n7270, B2 => n5099, C1 => n192, C2 => 
                           MEM_IN(23), A => n7368, ZN => n7367);
   U8042 : OAI22_X1 port map( A1 => n11318, A2 => n297, B1 => n5101, B2 => n144
                           , ZN => n7368);
   U8043 : AOI22_X1 port map( A1 => n7273, A2 => n5102, B1 => n7274, B2 => 
                           n5103, ZN => n7366);
   U8044 : AOI22_X1 port map( A1 => n7275, A2 => n5104, B1 => n7276, B2 => 
                           n5105, ZN => n7365);
   U8045 : NAND3_X1 port map( A1 => n7369, A2 => n7370, A3 => n7371, ZN => 
                           n12680);
   U8046 : AOI221_X1 port map( B1 => n7270, B2 => n5109, C1 => n192, C2 => 
                           MEM_IN(24), A => n7372, ZN => n7371);
   U8047 : OAI22_X1 port map( A1 => n11317, A2 => n297, B1 => n5111, B2 => n144
                           , ZN => n7372);
   U8048 : AOI22_X1 port map( A1 => n7273, A2 => n5112, B1 => n7274, B2 => 
                           n5113, ZN => n7370);
   U8049 : AOI22_X1 port map( A1 => n7275, A2 => n5114, B1 => n7276, B2 => 
                           n5115, ZN => n7369);
   U8050 : NAND3_X1 port map( A1 => n7373, A2 => n7374, A3 => n7375, ZN => 
                           n12679);
   U8051 : AOI221_X1 port map( B1 => n7270, B2 => n5119, C1 => n192, C2 => 
                           MEM_IN(25), A => n7376, ZN => n7375);
   U8052 : OAI22_X1 port map( A1 => n11316, A2 => n297, B1 => n5121, B2 => n144
                           , ZN => n7376);
   U8053 : AOI22_X1 port map( A1 => n7273, A2 => n5122, B1 => n7274, B2 => 
                           n5123, ZN => n7374);
   U8054 : AOI22_X1 port map( A1 => n7275, A2 => n5124, B1 => n7276, B2 => 
                           n5125, ZN => n7373);
   U8055 : NAND3_X1 port map( A1 => n7377, A2 => n7378, A3 => n7379, ZN => 
                           n12678);
   U8056 : AOI221_X1 port map( B1 => n7270, B2 => n5129, C1 => n192, C2 => 
                           MEM_IN(26), A => n7380, ZN => n7379);
   U8057 : OAI22_X1 port map( A1 => n11315, A2 => n297, B1 => n5131, B2 => n144
                           , ZN => n7380);
   U8058 : AOI22_X1 port map( A1 => n7273, A2 => n5132, B1 => n7274, B2 => 
                           n5133, ZN => n7378);
   U8059 : AOI22_X1 port map( A1 => n7275, A2 => n5134, B1 => n7276, B2 => 
                           n5135, ZN => n7377);
   U8060 : NAND3_X1 port map( A1 => n7381, A2 => n7382, A3 => n7383, ZN => 
                           n12677);
   U8061 : AOI221_X1 port map( B1 => n7270, B2 => n5139, C1 => n192, C2 => 
                           MEM_IN(27), A => n7384, ZN => n7383);
   U8062 : OAI22_X1 port map( A1 => n11314, A2 => n297, B1 => n5141, B2 => n144
                           , ZN => n7384);
   U8063 : AOI22_X1 port map( A1 => n7273, A2 => n5142, B1 => n7274, B2 => 
                           n5143, ZN => n7382);
   U8064 : AOI22_X1 port map( A1 => n7275, A2 => n5144, B1 => n7276, B2 => 
                           n5145, ZN => n7381);
   U8065 : NAND3_X1 port map( A1 => n7385, A2 => n7386, A3 => n7387, ZN => 
                           n12676);
   U8066 : AOI221_X1 port map( B1 => n7270, B2 => n5149, C1 => n192, C2 => 
                           MEM_IN(28), A => n7388, ZN => n7387);
   U8067 : OAI22_X1 port map( A1 => n11313, A2 => n297, B1 => n5151, B2 => n144
                           , ZN => n7388);
   U8068 : AOI22_X1 port map( A1 => n7273, A2 => n5152, B1 => n7274, B2 => 
                           n5153, ZN => n7386);
   U8069 : AOI22_X1 port map( A1 => n7275, A2 => n5154, B1 => n7276, B2 => 
                           n5155, ZN => n7385);
   U8070 : NAND3_X1 port map( A1 => n7389, A2 => n7390, A3 => n7391, ZN => 
                           n12675);
   U8071 : AOI221_X1 port map( B1 => n7270, B2 => n5159, C1 => n192, C2 => 
                           MEM_IN(29), A => n7392, ZN => n7391);
   U8072 : OAI22_X1 port map( A1 => n11312, A2 => n297, B1 => n5161, B2 => n144
                           , ZN => n7392);
   U8073 : AOI22_X1 port map( A1 => n7273, A2 => n5162, B1 => n7274, B2 => 
                           n5163, ZN => n7390);
   U8074 : AOI22_X1 port map( A1 => n7275, A2 => n5164, B1 => n7276, B2 => 
                           n5165, ZN => n7389);
   U8075 : NAND3_X1 port map( A1 => n7393, A2 => n7394, A3 => n7395, ZN => 
                           n12674);
   U8076 : AOI221_X1 port map( B1 => n7270, B2 => n5169, C1 => n192, C2 => 
                           MEM_IN(30), A => n7396, ZN => n7395);
   U8077 : OAI22_X1 port map( A1 => n11311, A2 => n297, B1 => n5171, B2 => n144
                           , ZN => n7396);
   U8078 : AOI22_X1 port map( A1 => n7273, A2 => n5172, B1 => n7274, B2 => 
                           n5173, ZN => n7394);
   U8079 : AOI22_X1 port map( A1 => n7275, A2 => n5174, B1 => n7276, B2 => 
                           n5175, ZN => n7393);
   U8080 : NAND3_X1 port map( A1 => n7397, A2 => n7398, A3 => n7399, ZN => 
                           n12673);
   U8081 : AOI221_X1 port map( B1 => n7270, B2 => n5179, C1 => n192, C2 => 
                           MEM_IN(31), A => n7400, ZN => n7399);
   U8082 : OAI22_X1 port map( A1 => n11310, A2 => n297, B1 => n5181, B2 => n144
                           , ZN => n7400);
   U8083 : INV_X1 port map( A => n7404, ZN => n7403);
   U8084 : INV_X1 port map( A => n6964, ZN => n6961);
   U8085 : AOI22_X1 port map( A1 => n7273, A2 => n5191, B1 => n7274, B2 => 
                           n5192, ZN => n7398);
   U8086 : AOI22_X1 port map( A1 => n7275, A2 => n5195, B1 => n7276, B2 => 
                           n5196, ZN => n7397);
   U8087 : OAI22_X1 port map( A1 => n7404, A2 => n7402, B1 => n208, B2 => n296,
                           ZN => n7405);
   U8088 : NAND3_X1 port map( A1 => n208, A2 => n297, A3 => n6379, ZN => n7402)
                           ;
   U8089 : INV_X1 port map( A => n7401, ZN => n6379);
   U8090 : OAI22_X1 port map( A1 => n4786, A2 => n7408, B1 => n7409, B2 => 
                           n5204, ZN => n7272);
   U8091 : NOR2_X1 port map( A1 => n7401, A2 => n7404, ZN => n7409);
   U8092 : NAND3_X1 port map( A1 => n7117, A2 => n6530, A3 => n7410, ZN => 
                           n7401);
   U8093 : AOI211_X1 port map( C1 => n6527, C2 => n6223, A => n7411, B => n6964
                           , ZN => n7408);
   U8094 : NAND2_X1 port map( A1 => n7412, A2 => n7413, ZN => n7404);
   U8095 : NOR2_X1 port map( A1 => n6530, A2 => n4787, ZN => n6964);
   U8096 : NAND2_X1 port map( A1 => n6228, A2 => n6531, ZN => n6530);
   U8097 : NAND3_X1 port map( A1 => n7414, A2 => n7415, A3 => n7416, ZN => 
                           n12672);
   U8098 : AOI221_X1 port map( B1 => n7417, B2 => n4863, C1 => n193, C2 => 
                           MEM_IN(0), A => n7418, ZN => n7416);
   U8099 : OAI22_X1 port map( A1 => n11309, A2 => n299, B1 => n4867, B2 => n145
                           , ZN => n7418);
   U8100 : AOI22_X1 port map( A1 => n7420, A2 => n4869, B1 => n7421, B2 => 
                           n4871, ZN => n7415);
   U8101 : AOI22_X1 port map( A1 => n7422, A2 => n4873, B1 => n7423, B2 => 
                           n4875, ZN => n7414);
   U8102 : NAND3_X1 port map( A1 => n7424, A2 => n7425, A3 => n7426, ZN => 
                           n12671);
   U8103 : AOI221_X1 port map( B1 => n7417, B2 => n4879, C1 => n193, C2 => 
                           MEM_IN(1), A => n7427, ZN => n7426);
   U8104 : OAI22_X1 port map( A1 => n11308, A2 => n299, B1 => n4881, B2 => n145
                           , ZN => n7427);
   U8105 : AOI22_X1 port map( A1 => n7420, A2 => n4882, B1 => n7421, B2 => 
                           n4883, ZN => n7425);
   U8106 : AOI22_X1 port map( A1 => n7422, A2 => n4884, B1 => n7423, B2 => 
                           n4885, ZN => n7424);
   U8107 : NAND3_X1 port map( A1 => n7428, A2 => n7429, A3 => n7430, ZN => 
                           n12670);
   U8108 : AOI221_X1 port map( B1 => n7417, B2 => n4889, C1 => n193, C2 => 
                           MEM_IN(2), A => n7431, ZN => n7430);
   U8109 : OAI22_X1 port map( A1 => n11307, A2 => n299, B1 => n4891, B2 => n145
                           , ZN => n7431);
   U8110 : AOI22_X1 port map( A1 => n7420, A2 => n4892, B1 => n7421, B2 => 
                           n4893, ZN => n7429);
   U8111 : AOI22_X1 port map( A1 => n7422, A2 => n4894, B1 => n7423, B2 => 
                           n4895, ZN => n7428);
   U8112 : NAND3_X1 port map( A1 => n7432, A2 => n7433, A3 => n7434, ZN => 
                           n12669);
   U8113 : AOI221_X1 port map( B1 => n7417, B2 => n4899, C1 => n193, C2 => 
                           MEM_IN(3), A => n7435, ZN => n7434);
   U8114 : OAI22_X1 port map( A1 => n11306, A2 => n299, B1 => n4901, B2 => n145
                           , ZN => n7435);
   U8115 : AOI22_X1 port map( A1 => n7420, A2 => n4902, B1 => n7421, B2 => 
                           n4903, ZN => n7433);
   U8116 : AOI22_X1 port map( A1 => n7422, A2 => n4904, B1 => n7423, B2 => 
                           n4905, ZN => n7432);
   U8117 : NAND3_X1 port map( A1 => n7436, A2 => n7437, A3 => n7438, ZN => 
                           n12668);
   U8118 : AOI221_X1 port map( B1 => n7417, B2 => n4909, C1 => n193, C2 => 
                           MEM_IN(4), A => n7439, ZN => n7438);
   U8119 : OAI22_X1 port map( A1 => n11305, A2 => n299, B1 => n4911, B2 => n145
                           , ZN => n7439);
   U8120 : AOI22_X1 port map( A1 => n7420, A2 => n4912, B1 => n7421, B2 => 
                           n4913, ZN => n7437);
   U8121 : AOI22_X1 port map( A1 => n7422, A2 => n4914, B1 => n7423, B2 => 
                           n4915, ZN => n7436);
   U8122 : NAND3_X1 port map( A1 => n7440, A2 => n7441, A3 => n7442, ZN => 
                           n12667);
   U8123 : AOI221_X1 port map( B1 => n7417, B2 => n4919, C1 => n193, C2 => 
                           MEM_IN(5), A => n7443, ZN => n7442);
   U8124 : OAI22_X1 port map( A1 => n11304, A2 => n299, B1 => n4921, B2 => n145
                           , ZN => n7443);
   U8125 : AOI22_X1 port map( A1 => n7420, A2 => n4922, B1 => n7421, B2 => 
                           n4923, ZN => n7441);
   U8126 : AOI22_X1 port map( A1 => n7422, A2 => n4924, B1 => n7423, B2 => 
                           n4925, ZN => n7440);
   U8127 : NAND3_X1 port map( A1 => n7444, A2 => n7445, A3 => n7446, ZN => 
                           n12666);
   U8128 : AOI221_X1 port map( B1 => n7417, B2 => n4929, C1 => n193, C2 => 
                           MEM_IN(6), A => n7447, ZN => n7446);
   U8129 : OAI22_X1 port map( A1 => n11303, A2 => n299, B1 => n4931, B2 => n145
                           , ZN => n7447);
   U8130 : AOI22_X1 port map( A1 => n7420, A2 => n4932, B1 => n7421, B2 => 
                           n4933, ZN => n7445);
   U8131 : AOI22_X1 port map( A1 => n7422, A2 => n4934, B1 => n7423, B2 => 
                           n4935, ZN => n7444);
   U8132 : NAND3_X1 port map( A1 => n7448, A2 => n7449, A3 => n7450, ZN => 
                           n12665);
   U8133 : AOI221_X1 port map( B1 => n7417, B2 => n4939, C1 => n193, C2 => 
                           MEM_IN(7), A => n7451, ZN => n7450);
   U8134 : OAI22_X1 port map( A1 => n11302, A2 => n299, B1 => n4941, B2 => n145
                           , ZN => n7451);
   U8135 : AOI22_X1 port map( A1 => n7420, A2 => n4942, B1 => n7421, B2 => 
                           n4943, ZN => n7449);
   U8136 : AOI22_X1 port map( A1 => n7422, A2 => n4944, B1 => n7423, B2 => 
                           n4945, ZN => n7448);
   U8137 : NAND3_X1 port map( A1 => n7452, A2 => n7453, A3 => n7454, ZN => 
                           n12664);
   U8138 : AOI221_X1 port map( B1 => n7417, B2 => n4949, C1 => n193, C2 => 
                           MEM_IN(8), A => n7455, ZN => n7454);
   U8139 : OAI22_X1 port map( A1 => n11301, A2 => n299, B1 => n4951, B2 => n145
                           , ZN => n7455);
   U8140 : AOI22_X1 port map( A1 => n7420, A2 => n4952, B1 => n7421, B2 => 
                           n4953, ZN => n7453);
   U8141 : AOI22_X1 port map( A1 => n7422, A2 => n4954, B1 => n7423, B2 => 
                           n4955, ZN => n7452);
   U8142 : NAND3_X1 port map( A1 => n7456, A2 => n7457, A3 => n7458, ZN => 
                           n12663);
   U8143 : AOI221_X1 port map( B1 => n7417, B2 => n4959, C1 => n193, C2 => 
                           MEM_IN(9), A => n7459, ZN => n7458);
   U8144 : OAI22_X1 port map( A1 => n11300, A2 => n299, B1 => n4961, B2 => n145
                           , ZN => n7459);
   U8145 : AOI22_X1 port map( A1 => n7420, A2 => n4962, B1 => n7421, B2 => 
                           n4963, ZN => n7457);
   U8146 : AOI22_X1 port map( A1 => n7422, A2 => n4964, B1 => n7423, B2 => 
                           n4965, ZN => n7456);
   U8147 : NAND3_X1 port map( A1 => n7460, A2 => n7461, A3 => n7462, ZN => 
                           n12662);
   U8148 : AOI221_X1 port map( B1 => n7417, B2 => n4969, C1 => n193, C2 => 
                           MEM_IN(10), A => n7463, ZN => n7462);
   U8149 : OAI22_X1 port map( A1 => n11299, A2 => n299, B1 => n4971, B2 => n145
                           , ZN => n7463);
   U8150 : AOI22_X1 port map( A1 => n7420, A2 => n4972, B1 => n7421, B2 => 
                           n4973, ZN => n7461);
   U8151 : AOI22_X1 port map( A1 => n7422, A2 => n4974, B1 => n7423, B2 => 
                           n4975, ZN => n7460);
   U8152 : NAND3_X1 port map( A1 => n7464, A2 => n7465, A3 => n7466, ZN => 
                           n12661);
   U8153 : AOI221_X1 port map( B1 => n7417, B2 => n4979, C1 => n193, C2 => 
                           MEM_IN(11), A => n7467, ZN => n7466);
   U8154 : OAI22_X1 port map( A1 => n11298, A2 => n299, B1 => n4981, B2 => n145
                           , ZN => n7467);
   U8155 : AOI22_X1 port map( A1 => n7420, A2 => n4982, B1 => n7421, B2 => 
                           n4983, ZN => n7465);
   U8156 : AOI22_X1 port map( A1 => n7422, A2 => n4984, B1 => n7423, B2 => 
                           n4985, ZN => n7464);
   U8157 : NAND3_X1 port map( A1 => n7468, A2 => n7469, A3 => n7470, ZN => 
                           n12660);
   U8158 : AOI221_X1 port map( B1 => n7417, B2 => n4989, C1 => n193, C2 => 
                           MEM_IN(12), A => n7471, ZN => n7470);
   U8159 : OAI22_X1 port map( A1 => n11297, A2 => n299, B1 => n4991, B2 => n145
                           , ZN => n7471);
   U8160 : AOI22_X1 port map( A1 => n7420, A2 => n4992, B1 => n7421, B2 => 
                           n4993, ZN => n7469);
   U8161 : AOI22_X1 port map( A1 => n7422, A2 => n4994, B1 => n7423, B2 => 
                           n4995, ZN => n7468);
   U8162 : NAND3_X1 port map( A1 => n7472, A2 => n7473, A3 => n7474, ZN => 
                           n12659);
   U8163 : AOI221_X1 port map( B1 => n7417, B2 => n4999, C1 => n193, C2 => 
                           MEM_IN(13), A => n7475, ZN => n7474);
   U8164 : OAI22_X1 port map( A1 => n11296, A2 => n299, B1 => n5001, B2 => n145
                           , ZN => n7475);
   U8165 : AOI22_X1 port map( A1 => n7420, A2 => n5002, B1 => n7421, B2 => 
                           n5003, ZN => n7473);
   U8166 : AOI22_X1 port map( A1 => n7422, A2 => n5004, B1 => n7423, B2 => 
                           n5005, ZN => n7472);
   U8167 : NAND3_X1 port map( A1 => n7476, A2 => n7477, A3 => n7478, ZN => 
                           n12658);
   U8168 : AOI221_X1 port map( B1 => n7417, B2 => n5009, C1 => n193, C2 => 
                           MEM_IN(14), A => n7479, ZN => n7478);
   U8169 : OAI22_X1 port map( A1 => n11295, A2 => n299, B1 => n5011, B2 => n145
                           , ZN => n7479);
   U8170 : AOI22_X1 port map( A1 => n7420, A2 => n5012, B1 => n7421, B2 => 
                           n5013, ZN => n7477);
   U8171 : AOI22_X1 port map( A1 => n7422, A2 => n5014, B1 => n7423, B2 => 
                           n5015, ZN => n7476);
   U8172 : NAND3_X1 port map( A1 => n7480, A2 => n7481, A3 => n7482, ZN => 
                           n12657);
   U8173 : AOI221_X1 port map( B1 => n7417, B2 => n5019, C1 => n193, C2 => 
                           MEM_IN(15), A => n7483, ZN => n7482);
   U8174 : OAI22_X1 port map( A1 => n11294, A2 => n299, B1 => n5021, B2 => n145
                           , ZN => n7483);
   U8175 : AOI22_X1 port map( A1 => n7420, A2 => n5022, B1 => n7421, B2 => 
                           n5023, ZN => n7481);
   U8176 : AOI22_X1 port map( A1 => n7422, A2 => n5024, B1 => n7423, B2 => 
                           n5025, ZN => n7480);
   U8177 : NAND3_X1 port map( A1 => n7484, A2 => n7485, A3 => n7486, ZN => 
                           n12656);
   U8178 : AOI221_X1 port map( B1 => n7417, B2 => n5029, C1 => n193, C2 => 
                           MEM_IN(16), A => n7487, ZN => n7486);
   U8179 : OAI22_X1 port map( A1 => n11293, A2 => n299, B1 => n5031, B2 => n145
                           , ZN => n7487);
   U8180 : AOI22_X1 port map( A1 => n7420, A2 => n5032, B1 => n7421, B2 => 
                           n5033, ZN => n7485);
   U8181 : AOI22_X1 port map( A1 => n7422, A2 => n5034, B1 => n7423, B2 => 
                           n5035, ZN => n7484);
   U8182 : NAND3_X1 port map( A1 => n7488, A2 => n7489, A3 => n7490, ZN => 
                           n12655);
   U8183 : AOI221_X1 port map( B1 => n7417, B2 => n5039, C1 => n193, C2 => 
                           MEM_IN(17), A => n7491, ZN => n7490);
   U8184 : OAI22_X1 port map( A1 => n11292, A2 => n299, B1 => n5041, B2 => n145
                           , ZN => n7491);
   U8185 : AOI22_X1 port map( A1 => n7420, A2 => n5042, B1 => n7421, B2 => 
                           n5043, ZN => n7489);
   U8186 : AOI22_X1 port map( A1 => n7422, A2 => n5044, B1 => n7423, B2 => 
                           n5045, ZN => n7488);
   U8187 : NAND3_X1 port map( A1 => n7492, A2 => n7493, A3 => n7494, ZN => 
                           n12654);
   U8188 : AOI221_X1 port map( B1 => n7417, B2 => n5049, C1 => n193, C2 => 
                           MEM_IN(18), A => n7495, ZN => n7494);
   U8189 : OAI22_X1 port map( A1 => n11291, A2 => n299, B1 => n5051, B2 => n145
                           , ZN => n7495);
   U8190 : AOI22_X1 port map( A1 => n7420, A2 => n5052, B1 => n7421, B2 => 
                           n5053, ZN => n7493);
   U8191 : AOI22_X1 port map( A1 => n7422, A2 => n5054, B1 => n7423, B2 => 
                           n5055, ZN => n7492);
   U8192 : NAND3_X1 port map( A1 => n7496, A2 => n7497, A3 => n7498, ZN => 
                           n12653);
   U8193 : AOI221_X1 port map( B1 => n7417, B2 => n5059, C1 => n193, C2 => 
                           MEM_IN(19), A => n7499, ZN => n7498);
   U8194 : OAI22_X1 port map( A1 => n11290, A2 => n299, B1 => n5061, B2 => n145
                           , ZN => n7499);
   U8195 : AOI22_X1 port map( A1 => n7420, A2 => n5062, B1 => n7421, B2 => 
                           n5063, ZN => n7497);
   U8196 : AOI22_X1 port map( A1 => n7422, A2 => n5064, B1 => n7423, B2 => 
                           n5065, ZN => n7496);
   U8197 : NAND3_X1 port map( A1 => n7500, A2 => n7501, A3 => n7502, ZN => 
                           n12652);
   U8198 : AOI221_X1 port map( B1 => n7417, B2 => n5069, C1 => n193, C2 => 
                           MEM_IN(20), A => n7503, ZN => n7502);
   U8199 : OAI22_X1 port map( A1 => n11289, A2 => n299, B1 => n5071, B2 => n145
                           , ZN => n7503);
   U8200 : AOI22_X1 port map( A1 => n7420, A2 => n5072, B1 => n7421, B2 => 
                           n5073, ZN => n7501);
   U8201 : AOI22_X1 port map( A1 => n7422, A2 => n5074, B1 => n7423, B2 => 
                           n5075, ZN => n7500);
   U8202 : NAND3_X1 port map( A1 => n7504, A2 => n7505, A3 => n7506, ZN => 
                           n12651);
   U8203 : AOI221_X1 port map( B1 => n7417, B2 => n5079, C1 => n193, C2 => 
                           MEM_IN(21), A => n7507, ZN => n7506);
   U8204 : OAI22_X1 port map( A1 => n11288, A2 => n299, B1 => n5081, B2 => n145
                           , ZN => n7507);
   U8205 : AOI22_X1 port map( A1 => n7420, A2 => n5082, B1 => n7421, B2 => 
                           n5083, ZN => n7505);
   U8206 : AOI22_X1 port map( A1 => n7422, A2 => n5084, B1 => n7423, B2 => 
                           n5085, ZN => n7504);
   U8207 : NAND3_X1 port map( A1 => n7508, A2 => n7509, A3 => n7510, ZN => 
                           n12650);
   U8208 : AOI221_X1 port map( B1 => n7417, B2 => n5089, C1 => n193, C2 => 
                           MEM_IN(22), A => n7511, ZN => n7510);
   U8209 : OAI22_X1 port map( A1 => n11287, A2 => n299, B1 => n5091, B2 => n145
                           , ZN => n7511);
   U8210 : AOI22_X1 port map( A1 => n7420, A2 => n5092, B1 => n7421, B2 => 
                           n5093, ZN => n7509);
   U8211 : AOI22_X1 port map( A1 => n7422, A2 => n5094, B1 => n7423, B2 => 
                           n5095, ZN => n7508);
   U8212 : NAND3_X1 port map( A1 => n7512, A2 => n7513, A3 => n7514, ZN => 
                           n12649);
   U8213 : AOI221_X1 port map( B1 => n7417, B2 => n5099, C1 => n193, C2 => 
                           MEM_IN(23), A => n7515, ZN => n7514);
   U8214 : OAI22_X1 port map( A1 => n11286, A2 => n299, B1 => n5101, B2 => n145
                           , ZN => n7515);
   U8215 : AOI22_X1 port map( A1 => n7420, A2 => n5102, B1 => n7421, B2 => 
                           n5103, ZN => n7513);
   U8216 : AOI22_X1 port map( A1 => n7422, A2 => n5104, B1 => n7423, B2 => 
                           n5105, ZN => n7512);
   U8217 : NAND3_X1 port map( A1 => n7516, A2 => n7517, A3 => n7518, ZN => 
                           n12648);
   U8218 : AOI221_X1 port map( B1 => n7417, B2 => n5109, C1 => n193, C2 => 
                           MEM_IN(24), A => n7519, ZN => n7518);
   U8219 : OAI22_X1 port map( A1 => n11285, A2 => n299, B1 => n5111, B2 => n145
                           , ZN => n7519);
   U8220 : AOI22_X1 port map( A1 => n7420, A2 => n5112, B1 => n7421, B2 => 
                           n5113, ZN => n7517);
   U8221 : AOI22_X1 port map( A1 => n7422, A2 => n5114, B1 => n7423, B2 => 
                           n5115, ZN => n7516);
   U8222 : NAND3_X1 port map( A1 => n7520, A2 => n7521, A3 => n7522, ZN => 
                           n12647);
   U8223 : AOI221_X1 port map( B1 => n7417, B2 => n5119, C1 => n193, C2 => 
                           MEM_IN(25), A => n7523, ZN => n7522);
   U8224 : OAI22_X1 port map( A1 => n11284, A2 => n299, B1 => n5121, B2 => n145
                           , ZN => n7523);
   U8225 : AOI22_X1 port map( A1 => n7420, A2 => n5122, B1 => n7421, B2 => 
                           n5123, ZN => n7521);
   U8226 : AOI22_X1 port map( A1 => n7422, A2 => n5124, B1 => n7423, B2 => 
                           n5125, ZN => n7520);
   U8227 : NAND3_X1 port map( A1 => n7524, A2 => n7525, A3 => n7526, ZN => 
                           n12646);
   U8228 : AOI221_X1 port map( B1 => n7417, B2 => n5129, C1 => n193, C2 => 
                           MEM_IN(26), A => n7527, ZN => n7526);
   U8229 : OAI22_X1 port map( A1 => n11283, A2 => n299, B1 => n5131, B2 => n145
                           , ZN => n7527);
   U8230 : AOI22_X1 port map( A1 => n7420, A2 => n5132, B1 => n7421, B2 => 
                           n5133, ZN => n7525);
   U8231 : AOI22_X1 port map( A1 => n7422, A2 => n5134, B1 => n7423, B2 => 
                           n5135, ZN => n7524);
   U8232 : NAND3_X1 port map( A1 => n7528, A2 => n7529, A3 => n7530, ZN => 
                           n12645);
   U8233 : AOI221_X1 port map( B1 => n7417, B2 => n5139, C1 => n193, C2 => 
                           MEM_IN(27), A => n7531, ZN => n7530);
   U8234 : OAI22_X1 port map( A1 => n11282, A2 => n299, B1 => n5141, B2 => n145
                           , ZN => n7531);
   U8235 : AOI22_X1 port map( A1 => n7420, A2 => n5142, B1 => n7421, B2 => 
                           n5143, ZN => n7529);
   U8236 : AOI22_X1 port map( A1 => n7422, A2 => n5144, B1 => n7423, B2 => 
                           n5145, ZN => n7528);
   U8237 : NAND3_X1 port map( A1 => n7532, A2 => n7533, A3 => n7534, ZN => 
                           n12644);
   U8238 : AOI221_X1 port map( B1 => n7417, B2 => n5149, C1 => n193, C2 => 
                           MEM_IN(28), A => n7535, ZN => n7534);
   U8239 : OAI22_X1 port map( A1 => n11281, A2 => n299, B1 => n5151, B2 => n145
                           , ZN => n7535);
   U8240 : AOI22_X1 port map( A1 => n7420, A2 => n5152, B1 => n7421, B2 => 
                           n5153, ZN => n7533);
   U8241 : AOI22_X1 port map( A1 => n7422, A2 => n5154, B1 => n7423, B2 => 
                           n5155, ZN => n7532);
   U8242 : NAND3_X1 port map( A1 => n7536, A2 => n7537, A3 => n7538, ZN => 
                           n12643);
   U8243 : AOI221_X1 port map( B1 => n7417, B2 => n5159, C1 => n193, C2 => 
                           MEM_IN(29), A => n7539, ZN => n7538);
   U8244 : OAI22_X1 port map( A1 => n11280, A2 => n299, B1 => n5161, B2 => n145
                           , ZN => n7539);
   U8245 : AOI22_X1 port map( A1 => n7420, A2 => n5162, B1 => n7421, B2 => 
                           n5163, ZN => n7537);
   U8246 : AOI22_X1 port map( A1 => n7422, A2 => n5164, B1 => n7423, B2 => 
                           n5165, ZN => n7536);
   U8247 : NAND3_X1 port map( A1 => n7540, A2 => n7541, A3 => n7542, ZN => 
                           n12642);
   U8248 : AOI221_X1 port map( B1 => n7417, B2 => n5169, C1 => n193, C2 => 
                           MEM_IN(30), A => n7543, ZN => n7542);
   U8249 : OAI22_X1 port map( A1 => n11279, A2 => n299, B1 => n5171, B2 => n145
                           , ZN => n7543);
   U8250 : AOI22_X1 port map( A1 => n7420, A2 => n5172, B1 => n7421, B2 => 
                           n5173, ZN => n7541);
   U8251 : AOI22_X1 port map( A1 => n7422, A2 => n5174, B1 => n7423, B2 => 
                           n5175, ZN => n7540);
   U8252 : NAND3_X1 port map( A1 => n7544, A2 => n7545, A3 => n7546, ZN => 
                           n12641);
   U8253 : AOI221_X1 port map( B1 => n7417, B2 => n5179, C1 => n193, C2 => 
                           MEM_IN(31), A => n7547, ZN => n7546);
   U8254 : OAI22_X1 port map( A1 => n11278, A2 => n299, B1 => n5181, B2 => n145
                           , ZN => n7547);
   U8255 : INV_X1 port map( A => n7551, ZN => n7550);
   U8256 : NAND2_X1 port map( A1 => n5206, A2 => n6969, ZN => n7260);
   U8257 : AOI22_X1 port map( A1 => n7420, A2 => n5191, B1 => n7421, B2 => 
                           n5192, ZN => n7545);
   U8258 : AOI22_X1 port map( A1 => n7422, A2 => n5195, B1 => n7423, B2 => 
                           n5196, ZN => n7544);
   U8259 : OAI22_X1 port map( A1 => n7551, A2 => n7549, B1 => n208, B2 => n298,
                           ZN => n7552);
   U8260 : NAND3_X1 port map( A1 => n208, A2 => n299, A3 => n6529, ZN => n7549)
                           ;
   U8261 : INV_X1 port map( A => n7548, ZN => n6529);
   U8262 : OAI22_X1 port map( A1 => n4786, A2 => n7555, B1 => n7556, B2 => 
                           n5204, ZN => n7419);
   U8263 : NOR2_X1 port map( A1 => n7548, A2 => n7551, ZN => n7556);
   U8264 : NAND2_X1 port map( A1 => n7557, A2 => n7117, ZN => n7548);
   U8265 : AOI211_X1 port map( C1 => n6527, C2 => n7558, A => n7411, B => n7554
                           , ZN => n7555);
   U8266 : OAI21_X1 port map( B1 => n7117, B2 => n4787, A => n5368, ZN => n7411
                           );
   U8267 : NOR2_X1 port map( A1 => n6969, A2 => n6973, ZN => n7117);
   U8268 : INV_X1 port map( A => n7559, ZN => n6973);
   U8269 : NAND2_X1 port map( A1 => n6823, A2 => n6678, ZN => n6969);
   U8270 : INV_X1 port map( A => n6971, ZN => n6527);
   U8271 : NAND3_X1 port map( A1 => n6378, A2 => n6377, A3 => n7560, ZN => 
                           n6971);
   U8272 : NAND2_X1 port map( A1 => n7561, A2 => n7562, ZN => n7551);
   U8273 : NOR2_X1 port map( A1 => n6678, A2 => n4787, ZN => n7113);
   U8274 : NAND2_X1 port map( A1 => n6381, A2 => n6531, ZN => n6678);
   U8275 : NAND3_X1 port map( A1 => n7563, A2 => n7564, A3 => n7565, ZN => 
                           n12640);
   U8276 : AOI221_X1 port map( B1 => n220, B2 => n4863, C1 => n186, C2 => 
                           MEM_IN(0), A => n7566, ZN => n7565);
   U8277 : OAI22_X1 port map( A1 => n11277, A2 => n263, B1 => n4867, B2 => n142
                           , ZN => n7566);
   U8278 : AOI22_X1 port map( A1 => n199, A2 => n4869, B1 => n161, B2 => n4871,
                           ZN => n7564);
   U8279 : AOI22_X1 port map( A1 => n241, A2 => n4873, B1 => n158, B2 => n4875,
                           ZN => n7563);
   U8280 : NAND3_X1 port map( A1 => n7568, A2 => n7569, A3 => n7570, ZN => 
                           n12639);
   U8281 : AOI221_X1 port map( B1 => n220, B2 => n4879, C1 => n186, C2 => 
                           MEM_IN(1), A => n7571, ZN => n7570);
   U8282 : OAI22_X1 port map( A1 => n11276, A2 => n263, B1 => n4881, B2 => n142
                           , ZN => n7571);
   U8283 : AOI22_X1 port map( A1 => n199, A2 => n4882, B1 => n161, B2 => n4883,
                           ZN => n7569);
   U8284 : AOI22_X1 port map( A1 => n241, A2 => n4884, B1 => n158, B2 => n4885,
                           ZN => n7568);
   U8285 : NAND3_X1 port map( A1 => n7572, A2 => n7573, A3 => n7574, ZN => 
                           n12638);
   U8286 : AOI221_X1 port map( B1 => n220, B2 => n4889, C1 => n186, C2 => 
                           MEM_IN(2), A => n7575, ZN => n7574);
   U8287 : OAI22_X1 port map( A1 => n11275, A2 => n263, B1 => n4891, B2 => n142
                           , ZN => n7575);
   U8288 : AOI22_X1 port map( A1 => n199, A2 => n4892, B1 => n161, B2 => n4893,
                           ZN => n7573);
   U8289 : AOI22_X1 port map( A1 => n241, A2 => n4894, B1 => n158, B2 => n4895,
                           ZN => n7572);
   U8290 : NAND3_X1 port map( A1 => n7576, A2 => n7577, A3 => n7578, ZN => 
                           n12637);
   U8291 : AOI221_X1 port map( B1 => n220, B2 => n4899, C1 => n186, C2 => 
                           MEM_IN(3), A => n7579, ZN => n7578);
   U8292 : OAI22_X1 port map( A1 => n11274, A2 => n263, B1 => n4901, B2 => n142
                           , ZN => n7579);
   U8293 : AOI22_X1 port map( A1 => n199, A2 => n4902, B1 => n161, B2 => n4903,
                           ZN => n7577);
   U8294 : AOI22_X1 port map( A1 => n241, A2 => n4904, B1 => n158, B2 => n4905,
                           ZN => n7576);
   U8295 : NAND3_X1 port map( A1 => n7580, A2 => n7581, A3 => n7582, ZN => 
                           n12636);
   U8296 : AOI221_X1 port map( B1 => n220, B2 => n4909, C1 => n186, C2 => 
                           MEM_IN(4), A => n7583, ZN => n7582);
   U8297 : OAI22_X1 port map( A1 => n11273, A2 => n263, B1 => n4911, B2 => n142
                           , ZN => n7583);
   U8298 : AOI22_X1 port map( A1 => n199, A2 => n4912, B1 => n161, B2 => n4913,
                           ZN => n7581);
   U8299 : AOI22_X1 port map( A1 => n241, A2 => n4914, B1 => n158, B2 => n4915,
                           ZN => n7580);
   U8300 : NAND3_X1 port map( A1 => n7584, A2 => n7585, A3 => n7586, ZN => 
                           n12635);
   U8301 : AOI221_X1 port map( B1 => n220, B2 => n4919, C1 => n186, C2 => 
                           MEM_IN(5), A => n7587, ZN => n7586);
   U8302 : OAI22_X1 port map( A1 => n11272, A2 => n263, B1 => n4921, B2 => n142
                           , ZN => n7587);
   U8303 : AOI22_X1 port map( A1 => n199, A2 => n4922, B1 => n161, B2 => n4923,
                           ZN => n7585);
   U8304 : AOI22_X1 port map( A1 => n241, A2 => n4924, B1 => n158, B2 => n4925,
                           ZN => n7584);
   U8305 : NAND3_X1 port map( A1 => n7588, A2 => n7589, A3 => n7590, ZN => 
                           n12634);
   U8306 : AOI221_X1 port map( B1 => n220, B2 => n4929, C1 => n186, C2 => 
                           MEM_IN(6), A => n7591, ZN => n7590);
   U8307 : OAI22_X1 port map( A1 => n11271, A2 => n263, B1 => n4931, B2 => n142
                           , ZN => n7591);
   U8308 : AOI22_X1 port map( A1 => n199, A2 => n4932, B1 => n161, B2 => n4933,
                           ZN => n7589);
   U8309 : AOI22_X1 port map( A1 => n241, A2 => n4934, B1 => n158, B2 => n4935,
                           ZN => n7588);
   U8310 : NAND3_X1 port map( A1 => n7592, A2 => n7593, A3 => n7594, ZN => 
                           n12633);
   U8311 : AOI221_X1 port map( B1 => n220, B2 => n4939, C1 => n186, C2 => 
                           MEM_IN(7), A => n7595, ZN => n7594);
   U8312 : OAI22_X1 port map( A1 => n11270, A2 => n263, B1 => n4941, B2 => n142
                           , ZN => n7595);
   U8313 : AOI22_X1 port map( A1 => n199, A2 => n4942, B1 => n161, B2 => n4943,
                           ZN => n7593);
   U8314 : AOI22_X1 port map( A1 => n241, A2 => n4944, B1 => n158, B2 => n4945,
                           ZN => n7592);
   U8315 : NAND3_X1 port map( A1 => n7596, A2 => n7597, A3 => n7598, ZN => 
                           n12632);
   U8316 : AOI221_X1 port map( B1 => n220, B2 => n4949, C1 => n186, C2 => 
                           MEM_IN(8), A => n7599, ZN => n7598);
   U8317 : OAI22_X1 port map( A1 => n11269, A2 => n263, B1 => n4951, B2 => n142
                           , ZN => n7599);
   U8318 : AOI22_X1 port map( A1 => n199, A2 => n4952, B1 => n161, B2 => n4953,
                           ZN => n7597);
   U8319 : AOI22_X1 port map( A1 => n241, A2 => n4954, B1 => n158, B2 => n4955,
                           ZN => n7596);
   U8320 : NAND3_X1 port map( A1 => n7600, A2 => n7601, A3 => n7602, ZN => 
                           n12631);
   U8321 : AOI221_X1 port map( B1 => n220, B2 => n4959, C1 => n186, C2 => 
                           MEM_IN(9), A => n7603, ZN => n7602);
   U8322 : OAI22_X1 port map( A1 => n11268, A2 => n263, B1 => n4961, B2 => n142
                           , ZN => n7603);
   U8323 : AOI22_X1 port map( A1 => n199, A2 => n4962, B1 => n161, B2 => n4963,
                           ZN => n7601);
   U8324 : AOI22_X1 port map( A1 => n241, A2 => n4964, B1 => n158, B2 => n4965,
                           ZN => n7600);
   U8325 : NAND3_X1 port map( A1 => n7604, A2 => n7605, A3 => n7606, ZN => 
                           n12630);
   U8326 : AOI221_X1 port map( B1 => n220, B2 => n4969, C1 => n186, C2 => 
                           MEM_IN(10), A => n7607, ZN => n7606);
   U8327 : OAI22_X1 port map( A1 => n11267, A2 => n263, B1 => n4971, B2 => n142
                           , ZN => n7607);
   U8328 : AOI22_X1 port map( A1 => n199, A2 => n4972, B1 => n161, B2 => n4973,
                           ZN => n7605);
   U8329 : AOI22_X1 port map( A1 => n241, A2 => n4974, B1 => n158, B2 => n4975,
                           ZN => n7604);
   U8330 : NAND3_X1 port map( A1 => n7608, A2 => n7609, A3 => n7610, ZN => 
                           n12629);
   U8331 : AOI221_X1 port map( B1 => n220, B2 => n4979, C1 => n186, C2 => 
                           MEM_IN(11), A => n7611, ZN => n7610);
   U8332 : OAI22_X1 port map( A1 => n11266, A2 => n263, B1 => n4981, B2 => n142
                           , ZN => n7611);
   U8333 : AOI22_X1 port map( A1 => n199, A2 => n4982, B1 => n161, B2 => n4983,
                           ZN => n7609);
   U8334 : AOI22_X1 port map( A1 => n241, A2 => n4984, B1 => n158, B2 => n4985,
                           ZN => n7608);
   U8335 : NAND3_X1 port map( A1 => n7612, A2 => n7613, A3 => n7614, ZN => 
                           n12628);
   U8336 : AOI221_X1 port map( B1 => n220, B2 => n4989, C1 => n186, C2 => 
                           MEM_IN(12), A => n7615, ZN => n7614);
   U8337 : OAI22_X1 port map( A1 => n11265, A2 => n263, B1 => n4991, B2 => n142
                           , ZN => n7615);
   U8338 : AOI22_X1 port map( A1 => n199, A2 => n4992, B1 => n161, B2 => n4993,
                           ZN => n7613);
   U8339 : AOI22_X1 port map( A1 => n241, A2 => n4994, B1 => n158, B2 => n4995,
                           ZN => n7612);
   U8340 : NAND3_X1 port map( A1 => n7616, A2 => n7617, A3 => n7618, ZN => 
                           n12627);
   U8341 : AOI221_X1 port map( B1 => n220, B2 => n4999, C1 => n186, C2 => 
                           MEM_IN(13), A => n7619, ZN => n7618);
   U8342 : OAI22_X1 port map( A1 => n11264, A2 => n263, B1 => n5001, B2 => n142
                           , ZN => n7619);
   U8343 : AOI22_X1 port map( A1 => n199, A2 => n5002, B1 => n161, B2 => n5003,
                           ZN => n7617);
   U8344 : AOI22_X1 port map( A1 => n241, A2 => n5004, B1 => n158, B2 => n5005,
                           ZN => n7616);
   U8345 : NAND3_X1 port map( A1 => n7620, A2 => n7621, A3 => n7622, ZN => 
                           n12626);
   U8346 : AOI221_X1 port map( B1 => n220, B2 => n5009, C1 => n186, C2 => 
                           MEM_IN(14), A => n7623, ZN => n7622);
   U8347 : OAI22_X1 port map( A1 => n11263, A2 => n263, B1 => n5011, B2 => n142
                           , ZN => n7623);
   U8348 : AOI22_X1 port map( A1 => n199, A2 => n5012, B1 => n161, B2 => n5013,
                           ZN => n7621);
   U8349 : AOI22_X1 port map( A1 => n241, A2 => n5014, B1 => n158, B2 => n5015,
                           ZN => n7620);
   U8350 : NAND3_X1 port map( A1 => n7624, A2 => n7625, A3 => n7626, ZN => 
                           n12625);
   U8351 : AOI221_X1 port map( B1 => n220, B2 => n5019, C1 => n186, C2 => 
                           MEM_IN(15), A => n7627, ZN => n7626);
   U8352 : OAI22_X1 port map( A1 => n11262, A2 => n263, B1 => n5021, B2 => n142
                           , ZN => n7627);
   U8353 : AOI22_X1 port map( A1 => n199, A2 => n5022, B1 => n161, B2 => n5023,
                           ZN => n7625);
   U8354 : AOI22_X1 port map( A1 => n241, A2 => n5024, B1 => n158, B2 => n5025,
                           ZN => n7624);
   U8355 : NAND3_X1 port map( A1 => n7628, A2 => n7629, A3 => n7630, ZN => 
                           n12624);
   U8356 : AOI221_X1 port map( B1 => n220, B2 => n5029, C1 => n186, C2 => 
                           MEM_IN(16), A => n7631, ZN => n7630);
   U8357 : OAI22_X1 port map( A1 => n11261, A2 => n263, B1 => n5031, B2 => n142
                           , ZN => n7631);
   U8358 : AOI22_X1 port map( A1 => n199, A2 => n5032, B1 => n161, B2 => n5033,
                           ZN => n7629);
   U8359 : AOI22_X1 port map( A1 => n241, A2 => n5034, B1 => n158, B2 => n5035,
                           ZN => n7628);
   U8360 : NAND3_X1 port map( A1 => n7632, A2 => n7633, A3 => n7634, ZN => 
                           n12623);
   U8361 : AOI221_X1 port map( B1 => n220, B2 => n5039, C1 => n186, C2 => 
                           MEM_IN(17), A => n7635, ZN => n7634);
   U8362 : OAI22_X1 port map( A1 => n11260, A2 => n263, B1 => n5041, B2 => n142
                           , ZN => n7635);
   U8363 : AOI22_X1 port map( A1 => n199, A2 => n5042, B1 => n161, B2 => n5043,
                           ZN => n7633);
   U8364 : AOI22_X1 port map( A1 => n241, A2 => n5044, B1 => n158, B2 => n5045,
                           ZN => n7632);
   U8365 : NAND3_X1 port map( A1 => n7636, A2 => n7637, A3 => n7638, ZN => 
                           n12622);
   U8366 : AOI221_X1 port map( B1 => n220, B2 => n5049, C1 => n186, C2 => 
                           MEM_IN(18), A => n7639, ZN => n7638);
   U8367 : OAI22_X1 port map( A1 => n11259, A2 => n263, B1 => n5051, B2 => n142
                           , ZN => n7639);
   U8368 : AOI22_X1 port map( A1 => n199, A2 => n5052, B1 => n161, B2 => n5053,
                           ZN => n7637);
   U8369 : AOI22_X1 port map( A1 => n241, A2 => n5054, B1 => n158, B2 => n5055,
                           ZN => n7636);
   U8370 : NAND3_X1 port map( A1 => n7640, A2 => n7641, A3 => n7642, ZN => 
                           n12621);
   U8371 : AOI221_X1 port map( B1 => n220, B2 => n5059, C1 => n186, C2 => 
                           MEM_IN(19), A => n7643, ZN => n7642);
   U8372 : OAI22_X1 port map( A1 => n11258, A2 => n263, B1 => n5061, B2 => n142
                           , ZN => n7643);
   U8373 : AOI22_X1 port map( A1 => n199, A2 => n5062, B1 => n161, B2 => n5063,
                           ZN => n7641);
   U8374 : AOI22_X1 port map( A1 => n241, A2 => n5064, B1 => n158, B2 => n5065,
                           ZN => n7640);
   U8375 : NAND3_X1 port map( A1 => n7644, A2 => n7645, A3 => n7646, ZN => 
                           n12620);
   U8376 : AOI221_X1 port map( B1 => n220, B2 => n5069, C1 => n186, C2 => 
                           MEM_IN(20), A => n7647, ZN => n7646);
   U8377 : OAI22_X1 port map( A1 => n11257, A2 => n263, B1 => n5071, B2 => n142
                           , ZN => n7647);
   U8378 : AOI22_X1 port map( A1 => n199, A2 => n5072, B1 => n161, B2 => n5073,
                           ZN => n7645);
   U8379 : AOI22_X1 port map( A1 => n241, A2 => n5074, B1 => n158, B2 => n5075,
                           ZN => n7644);
   U8380 : NAND3_X1 port map( A1 => n7648, A2 => n7649, A3 => n7650, ZN => 
                           n12619);
   U8381 : AOI221_X1 port map( B1 => n220, B2 => n5079, C1 => n186, C2 => 
                           MEM_IN(21), A => n7651, ZN => n7650);
   U8382 : OAI22_X1 port map( A1 => n11256, A2 => n263, B1 => n5081, B2 => n142
                           , ZN => n7651);
   U8383 : AOI22_X1 port map( A1 => n199, A2 => n5082, B1 => n161, B2 => n5083,
                           ZN => n7649);
   U8384 : AOI22_X1 port map( A1 => n241, A2 => n5084, B1 => n158, B2 => n5085,
                           ZN => n7648);
   U8385 : NAND3_X1 port map( A1 => n7652, A2 => n7653, A3 => n7654, ZN => 
                           n12618);
   U8386 : AOI221_X1 port map( B1 => n220, B2 => n5089, C1 => n186, C2 => 
                           MEM_IN(22), A => n7655, ZN => n7654);
   U8387 : OAI22_X1 port map( A1 => n11255, A2 => n263, B1 => n5091, B2 => n142
                           , ZN => n7655);
   U8388 : AOI22_X1 port map( A1 => n199, A2 => n5092, B1 => n161, B2 => n5093,
                           ZN => n7653);
   U8389 : AOI22_X1 port map( A1 => n241, A2 => n5094, B1 => n158, B2 => n5095,
                           ZN => n7652);
   U8390 : NAND3_X1 port map( A1 => n7656, A2 => n7657, A3 => n7658, ZN => 
                           n12617);
   U8391 : AOI221_X1 port map( B1 => n220, B2 => n5099, C1 => n186, C2 => 
                           MEM_IN(23), A => n7659, ZN => n7658);
   U8392 : OAI22_X1 port map( A1 => n11254, A2 => n263, B1 => n5101, B2 => n142
                           , ZN => n7659);
   U8393 : AOI22_X1 port map( A1 => n199, A2 => n5102, B1 => n161, B2 => n5103,
                           ZN => n7657);
   U8394 : AOI22_X1 port map( A1 => n241, A2 => n5104, B1 => n158, B2 => n5105,
                           ZN => n7656);
   U8395 : NAND3_X1 port map( A1 => n7660, A2 => n7661, A3 => n7662, ZN => 
                           n12616);
   U8396 : AOI221_X1 port map( B1 => n220, B2 => n5109, C1 => n186, C2 => 
                           MEM_IN(24), A => n7663, ZN => n7662);
   U8397 : OAI22_X1 port map( A1 => n11253, A2 => n263, B1 => n5111, B2 => n142
                           , ZN => n7663);
   U8398 : AOI22_X1 port map( A1 => n199, A2 => n5112, B1 => n161, B2 => n5113,
                           ZN => n7661);
   U8399 : AOI22_X1 port map( A1 => n241, A2 => n5114, B1 => n158, B2 => n5115,
                           ZN => n7660);
   U8400 : NAND3_X1 port map( A1 => n7664, A2 => n7665, A3 => n7666, ZN => 
                           n12615);
   U8401 : AOI221_X1 port map( B1 => n220, B2 => n5119, C1 => n186, C2 => 
                           MEM_IN(25), A => n7667, ZN => n7666);
   U8402 : OAI22_X1 port map( A1 => n11252, A2 => n263, B1 => n5121, B2 => n142
                           , ZN => n7667);
   U8403 : AOI22_X1 port map( A1 => n199, A2 => n5122, B1 => n161, B2 => n5123,
                           ZN => n7665);
   U8404 : AOI22_X1 port map( A1 => n241, A2 => n5124, B1 => n158, B2 => n5125,
                           ZN => n7664);
   U8405 : NAND3_X1 port map( A1 => n7668, A2 => n7669, A3 => n7670, ZN => 
                           n12614);
   U8406 : AOI221_X1 port map( B1 => n220, B2 => n5129, C1 => n186, C2 => 
                           MEM_IN(26), A => n7671, ZN => n7670);
   U8407 : OAI22_X1 port map( A1 => n11251, A2 => n263, B1 => n5131, B2 => n142
                           , ZN => n7671);
   U8408 : AOI22_X1 port map( A1 => n199, A2 => n5132, B1 => n161, B2 => n5133,
                           ZN => n7669);
   U8409 : AOI22_X1 port map( A1 => n241, A2 => n5134, B1 => n158, B2 => n5135,
                           ZN => n7668);
   U8410 : NAND3_X1 port map( A1 => n7672, A2 => n7673, A3 => n7674, ZN => 
                           n12613);
   U8411 : AOI221_X1 port map( B1 => n220, B2 => n5139, C1 => n186, C2 => 
                           MEM_IN(27), A => n7675, ZN => n7674);
   U8412 : OAI22_X1 port map( A1 => n11250, A2 => n263, B1 => n5141, B2 => n142
                           , ZN => n7675);
   U8413 : AOI22_X1 port map( A1 => n199, A2 => n5142, B1 => n161, B2 => n5143,
                           ZN => n7673);
   U8414 : AOI22_X1 port map( A1 => n241, A2 => n5144, B1 => n158, B2 => n5145,
                           ZN => n7672);
   U8415 : NAND3_X1 port map( A1 => n7676, A2 => n7677, A3 => n7678, ZN => 
                           n12612);
   U8416 : AOI221_X1 port map( B1 => n220, B2 => n5149, C1 => n186, C2 => 
                           MEM_IN(28), A => n7679, ZN => n7678);
   U8417 : OAI22_X1 port map( A1 => n11249, A2 => n263, B1 => n5151, B2 => n142
                           , ZN => n7679);
   U8418 : AOI22_X1 port map( A1 => n199, A2 => n5152, B1 => n161, B2 => n5153,
                           ZN => n7677);
   U8419 : AOI22_X1 port map( A1 => n241, A2 => n5154, B1 => n158, B2 => n5155,
                           ZN => n7676);
   U8420 : NAND3_X1 port map( A1 => n7680, A2 => n7681, A3 => n7682, ZN => 
                           n12611);
   U8421 : AOI221_X1 port map( B1 => n220, B2 => n5159, C1 => n186, C2 => 
                           MEM_IN(29), A => n7683, ZN => n7682);
   U8422 : OAI22_X1 port map( A1 => n11248, A2 => n263, B1 => n5161, B2 => n142
                           , ZN => n7683);
   U8423 : AOI22_X1 port map( A1 => n199, A2 => n5162, B1 => n161, B2 => n5163,
                           ZN => n7681);
   U8424 : AOI22_X1 port map( A1 => n241, A2 => n5164, B1 => n158, B2 => n5165,
                           ZN => n7680);
   U8425 : NAND3_X1 port map( A1 => n7684, A2 => n7685, A3 => n7686, ZN => 
                           n12610);
   U8426 : AOI221_X1 port map( B1 => n220, B2 => n5169, C1 => n186, C2 => 
                           MEM_IN(30), A => n7687, ZN => n7686);
   U8427 : OAI22_X1 port map( A1 => n11247, A2 => n263, B1 => n5171, B2 => n142
                           , ZN => n7687);
   U8428 : AOI22_X1 port map( A1 => n199, A2 => n5172, B1 => n161, B2 => n5173,
                           ZN => n7685);
   U8429 : AOI22_X1 port map( A1 => n241, A2 => n5174, B1 => n158, B2 => n5175,
                           ZN => n7684);
   U8430 : NAND3_X1 port map( A1 => n7688, A2 => n7689, A3 => n7690, ZN => 
                           n12609);
   U8431 : AOI221_X1 port map( B1 => n220, B2 => n5179, C1 => n186, C2 => 
                           MEM_IN(31), A => n7691, ZN => n7690);
   U8432 : OAI22_X1 port map( A1 => n11246, A2 => n263, B1 => n5181, B2 => n142
                           , ZN => n7691);
   U8433 : INV_X1 port map( A => n7697, ZN => n7696);
   U8434 : AOI22_X1 port map( A1 => n199, A2 => n5191, B1 => n161, B2 => n5192,
                           ZN => n7689);
   U8435 : AOI22_X1 port map( A1 => n241, A2 => n5195, B1 => n158, B2 => n5196,
                           ZN => n7688);
   U8436 : INV_X1 port map( A => n7407, ZN => n7406);
   U8437 : AOI22_X1 port map( A1 => n7694, A2 => n7700, B1 => n4841, B2 => n263
                           , ZN => n7695);
   U8438 : INV_X1 port map( A => n7693, ZN => n7700);
   U8439 : NAND3_X1 port map( A1 => n208, A2 => n263, A3 => n6677, ZN => n7693)
                           ;
   U8440 : INV_X1 port map( A => n7692, ZN => n6677);
   U8441 : OAI22_X1 port map( A1 => n4786, A2 => n7701, B1 => n7702, B2 => 
                           n5204, ZN => n7567);
   U8442 : NOR2_X1 port map( A1 => n7692, A2 => n7703, ZN => n7702);
   U8443 : NAND4_X1 port map( A1 => n7557, A2 => n7562, A3 => n7559, A4 => 
                           n6823, ZN => n7692);
   U8444 : AND4_X1 port map( A1 => n7704, A2 => n7553, A3 => n5368, A4 => n7698
                           , ZN => n7701);
   U8445 : INV_X1 port map( A => n7554, ZN => n7553);
   U8446 : AOI211_X1 port map( C1 => n5207, C2 => n7705, A => n7261, B => n7407
                           , ZN => n7704);
   U8447 : NOR2_X1 port map( A1 => n6823, A2 => n4787, ZN => n7261);
   U8448 : INV_X1 port map( A => n7703, ZN => n7694);
   U8449 : NAND2_X1 port map( A1 => n7706, A2 => n7707, ZN => n7703);
   U8450 : NAND2_X1 port map( A1 => n7708, A2 => n5215, ZN => n6823);
   U8451 : NAND3_X1 port map( A1 => n7709, A2 => n7710, A3 => n7711, ZN => 
                           n12608);
   U8452 : AOI221_X1 port map( B1 => n7712, B2 => n4863, C1 => n187, C2 => 
                           MEM_IN(0), A => n7713, ZN => n7711);
   U8453 : OAI22_X1 port map( A1 => n11245, A2 => n285, B1 => n4867, B2 => n143
                           , ZN => n7713);
   U8454 : AOI22_X1 port map( A1 => n7715, A2 => n4869, B1 => n7716, B2 => 
                           n4871, ZN => n7710);
   U8455 : AOI22_X1 port map( A1 => n7717, A2 => n4873, B1 => n7718, B2 => 
                           n4875, ZN => n7709);
   U8456 : NAND3_X1 port map( A1 => n7719, A2 => n7720, A3 => n7721, ZN => 
                           n12607);
   U8457 : AOI221_X1 port map( B1 => n7712, B2 => n4879, C1 => n187, C2 => 
                           MEM_IN(1), A => n7722, ZN => n7721);
   U8458 : OAI22_X1 port map( A1 => n11244, A2 => n285, B1 => n4881, B2 => n143
                           , ZN => n7722);
   U8459 : AOI22_X1 port map( A1 => n7715, A2 => n4882, B1 => n7716, B2 => 
                           n4883, ZN => n7720);
   U8460 : AOI22_X1 port map( A1 => n7717, A2 => n4884, B1 => n7718, B2 => 
                           n4885, ZN => n7719);
   U8461 : NAND3_X1 port map( A1 => n7723, A2 => n7724, A3 => n7725, ZN => 
                           n12606);
   U8462 : AOI221_X1 port map( B1 => n7712, B2 => n4889, C1 => n187, C2 => 
                           MEM_IN(2), A => n7726, ZN => n7725);
   U8463 : OAI22_X1 port map( A1 => n11243, A2 => n285, B1 => n4891, B2 => n143
                           , ZN => n7726);
   U8464 : AOI22_X1 port map( A1 => n7715, A2 => n4892, B1 => n7716, B2 => 
                           n4893, ZN => n7724);
   U8465 : AOI22_X1 port map( A1 => n7717, A2 => n4894, B1 => n7718, B2 => 
                           n4895, ZN => n7723);
   U8466 : NAND3_X1 port map( A1 => n7727, A2 => n7728, A3 => n7729, ZN => 
                           n12605);
   U8467 : AOI221_X1 port map( B1 => n7712, B2 => n4899, C1 => n187, C2 => 
                           MEM_IN(3), A => n7730, ZN => n7729);
   U8468 : OAI22_X1 port map( A1 => n11242, A2 => n285, B1 => n4901, B2 => n143
                           , ZN => n7730);
   U8469 : AOI22_X1 port map( A1 => n7715, A2 => n4902, B1 => n7716, B2 => 
                           n4903, ZN => n7728);
   U8470 : AOI22_X1 port map( A1 => n7717, A2 => n4904, B1 => n7718, B2 => 
                           n4905, ZN => n7727);
   U8471 : NAND3_X1 port map( A1 => n7731, A2 => n7732, A3 => n7733, ZN => 
                           n12604);
   U8472 : AOI221_X1 port map( B1 => n7712, B2 => n4909, C1 => n187, C2 => 
                           MEM_IN(4), A => n7734, ZN => n7733);
   U8473 : OAI22_X1 port map( A1 => n11241, A2 => n285, B1 => n4911, B2 => n143
                           , ZN => n7734);
   U8474 : AOI22_X1 port map( A1 => n7715, A2 => n4912, B1 => n7716, B2 => 
                           n4913, ZN => n7732);
   U8475 : AOI22_X1 port map( A1 => n7717, A2 => n4914, B1 => n7718, B2 => 
                           n4915, ZN => n7731);
   U8476 : NAND3_X1 port map( A1 => n7735, A2 => n7736, A3 => n7737, ZN => 
                           n12603);
   U8477 : AOI221_X1 port map( B1 => n7712, B2 => n4919, C1 => n187, C2 => 
                           MEM_IN(5), A => n7738, ZN => n7737);
   U8478 : OAI22_X1 port map( A1 => n11240, A2 => n285, B1 => n4921, B2 => n143
                           , ZN => n7738);
   U8479 : AOI22_X1 port map( A1 => n7715, A2 => n4922, B1 => n7716, B2 => 
                           n4923, ZN => n7736);
   U8480 : AOI22_X1 port map( A1 => n7717, A2 => n4924, B1 => n7718, B2 => 
                           n4925, ZN => n7735);
   U8481 : NAND3_X1 port map( A1 => n7739, A2 => n7740, A3 => n7741, ZN => 
                           n12602);
   U8482 : AOI221_X1 port map( B1 => n7712, B2 => n4929, C1 => n187, C2 => 
                           MEM_IN(6), A => n7742, ZN => n7741);
   U8483 : OAI22_X1 port map( A1 => n11239, A2 => n285, B1 => n4931, B2 => n143
                           , ZN => n7742);
   U8484 : AOI22_X1 port map( A1 => n7715, A2 => n4932, B1 => n7716, B2 => 
                           n4933, ZN => n7740);
   U8485 : AOI22_X1 port map( A1 => n7717, A2 => n4934, B1 => n7718, B2 => 
                           n4935, ZN => n7739);
   U8486 : NAND3_X1 port map( A1 => n7743, A2 => n7744, A3 => n7745, ZN => 
                           n12601);
   U8487 : AOI221_X1 port map( B1 => n7712, B2 => n4939, C1 => n187, C2 => 
                           MEM_IN(7), A => n7746, ZN => n7745);
   U8488 : OAI22_X1 port map( A1 => n11238, A2 => n285, B1 => n4941, B2 => n143
                           , ZN => n7746);
   U8489 : AOI22_X1 port map( A1 => n7715, A2 => n4942, B1 => n7716, B2 => 
                           n4943, ZN => n7744);
   U8490 : AOI22_X1 port map( A1 => n7717, A2 => n4944, B1 => n7718, B2 => 
                           n4945, ZN => n7743);
   U8491 : NAND3_X1 port map( A1 => n7747, A2 => n7748, A3 => n7749, ZN => 
                           n12600);
   U8492 : AOI221_X1 port map( B1 => n7712, B2 => n4949, C1 => n187, C2 => 
                           MEM_IN(8), A => n7750, ZN => n7749);
   U8493 : OAI22_X1 port map( A1 => n11237, A2 => n285, B1 => n4951, B2 => n143
                           , ZN => n7750);
   U8494 : AOI22_X1 port map( A1 => n7715, A2 => n4952, B1 => n7716, B2 => 
                           n4953, ZN => n7748);
   U8495 : AOI22_X1 port map( A1 => n7717, A2 => n4954, B1 => n7718, B2 => 
                           n4955, ZN => n7747);
   U8496 : NAND3_X1 port map( A1 => n7751, A2 => n7752, A3 => n7753, ZN => 
                           n12599);
   U8497 : AOI221_X1 port map( B1 => n7712, B2 => n4959, C1 => n187, C2 => 
                           MEM_IN(9), A => n7754, ZN => n7753);
   U8498 : OAI22_X1 port map( A1 => n11236, A2 => n285, B1 => n4961, B2 => n143
                           , ZN => n7754);
   U8499 : AOI22_X1 port map( A1 => n7715, A2 => n4962, B1 => n7716, B2 => 
                           n4963, ZN => n7752);
   U8500 : AOI22_X1 port map( A1 => n7717, A2 => n4964, B1 => n7718, B2 => 
                           n4965, ZN => n7751);
   U8501 : NAND3_X1 port map( A1 => n7755, A2 => n7756, A3 => n7757, ZN => 
                           n12598);
   U8502 : AOI221_X1 port map( B1 => n7712, B2 => n4969, C1 => n187, C2 => 
                           MEM_IN(10), A => n7758, ZN => n7757);
   U8503 : OAI22_X1 port map( A1 => n11235, A2 => n285, B1 => n4971, B2 => n143
                           , ZN => n7758);
   U8504 : AOI22_X1 port map( A1 => n7715, A2 => n4972, B1 => n7716, B2 => 
                           n4973, ZN => n7756);
   U8505 : AOI22_X1 port map( A1 => n7717, A2 => n4974, B1 => n7718, B2 => 
                           n4975, ZN => n7755);
   U8506 : NAND3_X1 port map( A1 => n7759, A2 => n7760, A3 => n7761, ZN => 
                           n12597);
   U8507 : AOI221_X1 port map( B1 => n7712, B2 => n4979, C1 => n187, C2 => 
                           MEM_IN(11), A => n7762, ZN => n7761);
   U8508 : OAI22_X1 port map( A1 => n11234, A2 => n285, B1 => n4981, B2 => n143
                           , ZN => n7762);
   U8509 : AOI22_X1 port map( A1 => n7715, A2 => n4982, B1 => n7716, B2 => 
                           n4983, ZN => n7760);
   U8510 : AOI22_X1 port map( A1 => n7717, A2 => n4984, B1 => n7718, B2 => 
                           n4985, ZN => n7759);
   U8511 : NAND3_X1 port map( A1 => n7763, A2 => n7764, A3 => n7765, ZN => 
                           n12596);
   U8512 : AOI221_X1 port map( B1 => n7712, B2 => n4989, C1 => n187, C2 => 
                           MEM_IN(12), A => n7766, ZN => n7765);
   U8513 : OAI22_X1 port map( A1 => n11233, A2 => n285, B1 => n4991, B2 => n143
                           , ZN => n7766);
   U8514 : AOI22_X1 port map( A1 => n7715, A2 => n4992, B1 => n7716, B2 => 
                           n4993, ZN => n7764);
   U8515 : AOI22_X1 port map( A1 => n7717, A2 => n4994, B1 => n7718, B2 => 
                           n4995, ZN => n7763);
   U8516 : NAND3_X1 port map( A1 => n7767, A2 => n7768, A3 => n7769, ZN => 
                           n12595);
   U8517 : AOI221_X1 port map( B1 => n7712, B2 => n4999, C1 => n187, C2 => 
                           MEM_IN(13), A => n7770, ZN => n7769);
   U8518 : OAI22_X1 port map( A1 => n11232, A2 => n285, B1 => n5001, B2 => n143
                           , ZN => n7770);
   U8519 : AOI22_X1 port map( A1 => n7715, A2 => n5002, B1 => n7716, B2 => 
                           n5003, ZN => n7768);
   U8520 : AOI22_X1 port map( A1 => n7717, A2 => n5004, B1 => n7718, B2 => 
                           n5005, ZN => n7767);
   U8521 : NAND3_X1 port map( A1 => n7771, A2 => n7772, A3 => n7773, ZN => 
                           n12594);
   U8522 : AOI221_X1 port map( B1 => n7712, B2 => n5009, C1 => n187, C2 => 
                           MEM_IN(14), A => n7774, ZN => n7773);
   U8523 : OAI22_X1 port map( A1 => n11231, A2 => n285, B1 => n5011, B2 => n143
                           , ZN => n7774);
   U8524 : AOI22_X1 port map( A1 => n7715, A2 => n5012, B1 => n7716, B2 => 
                           n5013, ZN => n7772);
   U8525 : AOI22_X1 port map( A1 => n7717, A2 => n5014, B1 => n7718, B2 => 
                           n5015, ZN => n7771);
   U8526 : NAND3_X1 port map( A1 => n7775, A2 => n7776, A3 => n7777, ZN => 
                           n12593);
   U8527 : AOI221_X1 port map( B1 => n7712, B2 => n5019, C1 => n187, C2 => 
                           MEM_IN(15), A => n7778, ZN => n7777);
   U8528 : OAI22_X1 port map( A1 => n11230, A2 => n285, B1 => n5021, B2 => n143
                           , ZN => n7778);
   U8529 : AOI22_X1 port map( A1 => n7715, A2 => n5022, B1 => n7716, B2 => 
                           n5023, ZN => n7776);
   U8530 : AOI22_X1 port map( A1 => n7717, A2 => n5024, B1 => n7718, B2 => 
                           n5025, ZN => n7775);
   U8531 : NAND3_X1 port map( A1 => n7779, A2 => n7780, A3 => n7781, ZN => 
                           n12592);
   U8532 : AOI221_X1 port map( B1 => n7712, B2 => n5029, C1 => n187, C2 => 
                           MEM_IN(16), A => n7782, ZN => n7781);
   U8533 : OAI22_X1 port map( A1 => n11229, A2 => n285, B1 => n5031, B2 => n143
                           , ZN => n7782);
   U8534 : AOI22_X1 port map( A1 => n7715, A2 => n5032, B1 => n7716, B2 => 
                           n5033, ZN => n7780);
   U8535 : AOI22_X1 port map( A1 => n7717, A2 => n5034, B1 => n7718, B2 => 
                           n5035, ZN => n7779);
   U8536 : NAND3_X1 port map( A1 => n7783, A2 => n7784, A3 => n7785, ZN => 
                           n12591);
   U8537 : AOI221_X1 port map( B1 => n7712, B2 => n5039, C1 => n187, C2 => 
                           MEM_IN(17), A => n7786, ZN => n7785);
   U8538 : OAI22_X1 port map( A1 => n11228, A2 => n285, B1 => n5041, B2 => n143
                           , ZN => n7786);
   U8539 : AOI22_X1 port map( A1 => n7715, A2 => n5042, B1 => n7716, B2 => 
                           n5043, ZN => n7784);
   U8540 : AOI22_X1 port map( A1 => n7717, A2 => n5044, B1 => n7718, B2 => 
                           n5045, ZN => n7783);
   U8541 : NAND3_X1 port map( A1 => n7787, A2 => n7788, A3 => n7789, ZN => 
                           n12590);
   U8542 : AOI221_X1 port map( B1 => n7712, B2 => n5049, C1 => n187, C2 => 
                           MEM_IN(18), A => n7790, ZN => n7789);
   U8543 : OAI22_X1 port map( A1 => n11227, A2 => n285, B1 => n5051, B2 => n143
                           , ZN => n7790);
   U8544 : AOI22_X1 port map( A1 => n7715, A2 => n5052, B1 => n7716, B2 => 
                           n5053, ZN => n7788);
   U8545 : AOI22_X1 port map( A1 => n7717, A2 => n5054, B1 => n7718, B2 => 
                           n5055, ZN => n7787);
   U8546 : NAND3_X1 port map( A1 => n7791, A2 => n7792, A3 => n7793, ZN => 
                           n12589);
   U8547 : AOI221_X1 port map( B1 => n7712, B2 => n5059, C1 => n187, C2 => 
                           MEM_IN(19), A => n7794, ZN => n7793);
   U8548 : OAI22_X1 port map( A1 => n11226, A2 => n285, B1 => n5061, B2 => n143
                           , ZN => n7794);
   U8549 : AOI22_X1 port map( A1 => n7715, A2 => n5062, B1 => n7716, B2 => 
                           n5063, ZN => n7792);
   U8550 : AOI22_X1 port map( A1 => n7717, A2 => n5064, B1 => n7718, B2 => 
                           n5065, ZN => n7791);
   U8551 : NAND3_X1 port map( A1 => n7795, A2 => n7796, A3 => n7797, ZN => 
                           n12588);
   U8552 : AOI221_X1 port map( B1 => n7712, B2 => n5069, C1 => n187, C2 => 
                           MEM_IN(20), A => n7798, ZN => n7797);
   U8553 : OAI22_X1 port map( A1 => n11225, A2 => n285, B1 => n5071, B2 => n143
                           , ZN => n7798);
   U8554 : AOI22_X1 port map( A1 => n7715, A2 => n5072, B1 => n7716, B2 => 
                           n5073, ZN => n7796);
   U8555 : AOI22_X1 port map( A1 => n7717, A2 => n5074, B1 => n7718, B2 => 
                           n5075, ZN => n7795);
   U8556 : NAND3_X1 port map( A1 => n7799, A2 => n7800, A3 => n7801, ZN => 
                           n12587);
   U8557 : AOI221_X1 port map( B1 => n7712, B2 => n5079, C1 => n187, C2 => 
                           MEM_IN(21), A => n7802, ZN => n7801);
   U8558 : OAI22_X1 port map( A1 => n11224, A2 => n285, B1 => n5081, B2 => n143
                           , ZN => n7802);
   U8559 : AOI22_X1 port map( A1 => n7715, A2 => n5082, B1 => n7716, B2 => 
                           n5083, ZN => n7800);
   U8560 : AOI22_X1 port map( A1 => n7717, A2 => n5084, B1 => n7718, B2 => 
                           n5085, ZN => n7799);
   U8561 : NAND3_X1 port map( A1 => n7803, A2 => n7804, A3 => n7805, ZN => 
                           n12586);
   U8562 : AOI221_X1 port map( B1 => n7712, B2 => n5089, C1 => n187, C2 => 
                           MEM_IN(22), A => n7806, ZN => n7805);
   U8563 : OAI22_X1 port map( A1 => n11223, A2 => n285, B1 => n5091, B2 => n143
                           , ZN => n7806);
   U8564 : AOI22_X1 port map( A1 => n7715, A2 => n5092, B1 => n7716, B2 => 
                           n5093, ZN => n7804);
   U8565 : AOI22_X1 port map( A1 => n7717, A2 => n5094, B1 => n7718, B2 => 
                           n5095, ZN => n7803);
   U8566 : NAND3_X1 port map( A1 => n7807, A2 => n7808, A3 => n7809, ZN => 
                           n12585);
   U8567 : AOI221_X1 port map( B1 => n7712, B2 => n5099, C1 => n187, C2 => 
                           MEM_IN(23), A => n7810, ZN => n7809);
   U8568 : OAI22_X1 port map( A1 => n11222, A2 => n285, B1 => n5101, B2 => n143
                           , ZN => n7810);
   U8569 : AOI22_X1 port map( A1 => n7715, A2 => n5102, B1 => n7716, B2 => 
                           n5103, ZN => n7808);
   U8570 : AOI22_X1 port map( A1 => n7717, A2 => n5104, B1 => n7718, B2 => 
                           n5105, ZN => n7807);
   U8571 : NAND3_X1 port map( A1 => n7811, A2 => n7812, A3 => n7813, ZN => 
                           n12584);
   U8572 : AOI221_X1 port map( B1 => n7712, B2 => n5109, C1 => n187, C2 => 
                           MEM_IN(24), A => n7814, ZN => n7813);
   U8573 : OAI22_X1 port map( A1 => n11221, A2 => n285, B1 => n5111, B2 => n143
                           , ZN => n7814);
   U8574 : AOI22_X1 port map( A1 => n7715, A2 => n5112, B1 => n7716, B2 => 
                           n5113, ZN => n7812);
   U8575 : AOI22_X1 port map( A1 => n7717, A2 => n5114, B1 => n7718, B2 => 
                           n5115, ZN => n7811);
   U8576 : NAND3_X1 port map( A1 => n7815, A2 => n7816, A3 => n7817, ZN => 
                           n12583);
   U8577 : AOI221_X1 port map( B1 => n7712, B2 => n5119, C1 => n187, C2 => 
                           MEM_IN(25), A => n7818, ZN => n7817);
   U8578 : OAI22_X1 port map( A1 => n11220, A2 => n285, B1 => n5121, B2 => n143
                           , ZN => n7818);
   U8579 : AOI22_X1 port map( A1 => n7715, A2 => n5122, B1 => n7716, B2 => 
                           n5123, ZN => n7816);
   U8580 : AOI22_X1 port map( A1 => n7717, A2 => n5124, B1 => n7718, B2 => 
                           n5125, ZN => n7815);
   U8581 : NAND3_X1 port map( A1 => n7819, A2 => n7820, A3 => n7821, ZN => 
                           n12582);
   U8582 : AOI221_X1 port map( B1 => n7712, B2 => n5129, C1 => n187, C2 => 
                           MEM_IN(26), A => n7822, ZN => n7821);
   U8583 : OAI22_X1 port map( A1 => n11219, A2 => n285, B1 => n5131, B2 => n143
                           , ZN => n7822);
   U8584 : AOI22_X1 port map( A1 => n7715, A2 => n5132, B1 => n7716, B2 => 
                           n5133, ZN => n7820);
   U8585 : AOI22_X1 port map( A1 => n7717, A2 => n5134, B1 => n7718, B2 => 
                           n5135, ZN => n7819);
   U8586 : NAND3_X1 port map( A1 => n7823, A2 => n7824, A3 => n7825, ZN => 
                           n12581);
   U8587 : AOI221_X1 port map( B1 => n7712, B2 => n5139, C1 => n187, C2 => 
                           MEM_IN(27), A => n7826, ZN => n7825);
   U8588 : OAI22_X1 port map( A1 => n11218, A2 => n285, B1 => n5141, B2 => n143
                           , ZN => n7826);
   U8589 : AOI22_X1 port map( A1 => n7715, A2 => n5142, B1 => n7716, B2 => 
                           n5143, ZN => n7824);
   U8590 : AOI22_X1 port map( A1 => n7717, A2 => n5144, B1 => n7718, B2 => 
                           n5145, ZN => n7823);
   U8591 : NAND3_X1 port map( A1 => n7827, A2 => n7828, A3 => n7829, ZN => 
                           n12580);
   U8592 : AOI221_X1 port map( B1 => n7712, B2 => n5149, C1 => n187, C2 => 
                           MEM_IN(28), A => n7830, ZN => n7829);
   U8593 : OAI22_X1 port map( A1 => n11217, A2 => n285, B1 => n5151, B2 => n143
                           , ZN => n7830);
   U8594 : AOI22_X1 port map( A1 => n7715, A2 => n5152, B1 => n7716, B2 => 
                           n5153, ZN => n7828);
   U8595 : AOI22_X1 port map( A1 => n7717, A2 => n5154, B1 => n7718, B2 => 
                           n5155, ZN => n7827);
   U8596 : NAND3_X1 port map( A1 => n7831, A2 => n7832, A3 => n7833, ZN => 
                           n12579);
   U8597 : AOI221_X1 port map( B1 => n7712, B2 => n5159, C1 => n187, C2 => 
                           MEM_IN(29), A => n7834, ZN => n7833);
   U8598 : OAI22_X1 port map( A1 => n11216, A2 => n285, B1 => n5161, B2 => n143
                           , ZN => n7834);
   U8599 : AOI22_X1 port map( A1 => n7715, A2 => n5162, B1 => n7716, B2 => 
                           n5163, ZN => n7832);
   U8600 : AOI22_X1 port map( A1 => n7717, A2 => n5164, B1 => n7718, B2 => 
                           n5165, ZN => n7831);
   U8601 : NAND3_X1 port map( A1 => n7835, A2 => n7836, A3 => n7837, ZN => 
                           n12578);
   U8602 : AOI221_X1 port map( B1 => n7712, B2 => n5169, C1 => n187, C2 => 
                           MEM_IN(30), A => n7838, ZN => n7837);
   U8603 : OAI22_X1 port map( A1 => n11215, A2 => n285, B1 => n5171, B2 => n143
                           , ZN => n7838);
   U8604 : AOI22_X1 port map( A1 => n7715, A2 => n5172, B1 => n7716, B2 => 
                           n5173, ZN => n7836);
   U8605 : AOI22_X1 port map( A1 => n7717, A2 => n5174, B1 => n7718, B2 => 
                           n5175, ZN => n7835);
   U8606 : NAND3_X1 port map( A1 => n7839, A2 => n7840, A3 => n7841, ZN => 
                           n12577);
   U8607 : AOI221_X1 port map( B1 => n7712, B2 => n5179, C1 => n187, C2 => 
                           MEM_IN(31), A => n7842, ZN => n7841);
   U8608 : OAI22_X1 port map( A1 => n11214, A2 => n285, B1 => n5181, B2 => n143
                           , ZN => n7842);
   U8609 : INV_X1 port map( A => n7846, ZN => n7845);
   U8610 : NAND2_X1 port map( A1 => n5206, A2 => n7699, ZN => n7697);
   U8611 : NAND3_X1 port map( A1 => n5206, A2 => n7559, A3 => n7410, ZN => 
                           n7699);
   U8612 : AOI22_X1 port map( A1 => n7715, A2 => n5191, B1 => n7716, B2 => 
                           n5192, ZN => n7840);
   U8613 : AOI22_X1 port map( A1 => n7717, A2 => n5195, B1 => n7718, B2 => 
                           n5196, ZN => n7839);
   U8614 : OAI22_X1 port map( A1 => n7846, A2 => n7844, B1 => n208, B2 => n284,
                           ZN => n7848);
   U8615 : NAND3_X1 port map( A1 => n208, A2 => n285, A3 => n6822, ZN => n7844)
                           ;
   U8616 : INV_X1 port map( A => n7843, ZN => n6822);
   U8617 : OAI22_X1 port map( A1 => n4786, A2 => n7851, B1 => n7852, B2 => 
                           n5204, ZN => n7714);
   U8618 : NOR2_X1 port map( A1 => n7843, A2 => n7846, ZN => n7852);
   U8619 : NAND3_X1 port map( A1 => n7557, A2 => n7559, A3 => n7853, ZN => 
                           n7843);
   U8620 : NOR3_X1 port map( A1 => n7854, A2 => RESET, A3 => n7407, ZN => n7851
                           );
   U8621 : OAI22_X1 port map( A1 => n7855, A2 => n7856, B1 => n7557, B2 => 
                           n4787, ZN => n7854);
   U8622 : NAND2_X1 port map( A1 => n7857, A2 => n7858, ZN => n7846);
   U8623 : NOR2_X1 port map( A1 => n7559, A2 => n4787, ZN => n7407);
   U8624 : NAND2_X1 port map( A1 => n7708, A2 => n5372, ZN => n7559);
   U8625 : NAND3_X1 port map( A1 => n7859, A2 => n7860, A3 => n7861, ZN => 
                           n12576);
   U8626 : AOI221_X1 port map( B1 => n7862, B2 => n4863, C1 => n7863, C2 => 
                           MEM_IN(0), A => n7864, ZN => n7861);
   U8627 : OAI22_X1 port map( A1 => n11213, A2 => n218, B1 => n4867, B2 => n140
                           , ZN => n7864);
   U8628 : AOI22_X1 port map( A1 => n7866, A2 => n4869, B1 => n7867, B2 => 
                           n4871, ZN => n7860);
   U8629 : AOI22_X1 port map( A1 => n7868, A2 => n4873, B1 => n7869, B2 => 
                           n4875, ZN => n7859);
   U8630 : NAND3_X1 port map( A1 => n7870, A2 => n7871, A3 => n7872, ZN => 
                           n12575);
   U8631 : AOI221_X1 port map( B1 => n7862, B2 => n4879, C1 => n7863, C2 => 
                           MEM_IN(1), A => n7873, ZN => n7872);
   U8632 : OAI22_X1 port map( A1 => n11212, A2 => n218, B1 => n4881, B2 => n140
                           , ZN => n7873);
   U8633 : AOI22_X1 port map( A1 => n7866, A2 => n4882, B1 => n7867, B2 => 
                           n4883, ZN => n7871);
   U8634 : AOI22_X1 port map( A1 => n7868, A2 => n4884, B1 => n7869, B2 => 
                           n4885, ZN => n7870);
   U8635 : NAND3_X1 port map( A1 => n7874, A2 => n7875, A3 => n7876, ZN => 
                           n12574);
   U8636 : AOI221_X1 port map( B1 => n7862, B2 => n4889, C1 => n7863, C2 => 
                           MEM_IN(2), A => n7877, ZN => n7876);
   U8637 : OAI22_X1 port map( A1 => n11211, A2 => n218, B1 => n4891, B2 => n140
                           , ZN => n7877);
   U8638 : AOI22_X1 port map( A1 => n7866, A2 => n4892, B1 => n7867, B2 => 
                           n4893, ZN => n7875);
   U8639 : AOI22_X1 port map( A1 => n7868, A2 => n4894, B1 => n7869, B2 => 
                           n4895, ZN => n7874);
   U8640 : NAND3_X1 port map( A1 => n7878, A2 => n7879, A3 => n7880, ZN => 
                           n12573);
   U8641 : AOI221_X1 port map( B1 => n7862, B2 => n4899, C1 => n7863, C2 => 
                           MEM_IN(3), A => n7881, ZN => n7880);
   U8642 : OAI22_X1 port map( A1 => n11210, A2 => n218, B1 => n4901, B2 => n140
                           , ZN => n7881);
   U8643 : AOI22_X1 port map( A1 => n7866, A2 => n4902, B1 => n7867, B2 => 
                           n4903, ZN => n7879);
   U8644 : AOI22_X1 port map( A1 => n7868, A2 => n4904, B1 => n7869, B2 => 
                           n4905, ZN => n7878);
   U8645 : NAND3_X1 port map( A1 => n7882, A2 => n7883, A3 => n7884, ZN => 
                           n12572);
   U8646 : AOI221_X1 port map( B1 => n7862, B2 => n4909, C1 => n7863, C2 => 
                           MEM_IN(4), A => n7885, ZN => n7884);
   U8647 : OAI22_X1 port map( A1 => n11209, A2 => n218, B1 => n4911, B2 => n140
                           , ZN => n7885);
   U8648 : AOI22_X1 port map( A1 => n7866, A2 => n4912, B1 => n7867, B2 => 
                           n4913, ZN => n7883);
   U8649 : AOI22_X1 port map( A1 => n7868, A2 => n4914, B1 => n7869, B2 => 
                           n4915, ZN => n7882);
   U8650 : NAND3_X1 port map( A1 => n7886, A2 => n7887, A3 => n7888, ZN => 
                           n12571);
   U8651 : AOI221_X1 port map( B1 => n7862, B2 => n4919, C1 => n7863, C2 => 
                           MEM_IN(5), A => n7889, ZN => n7888);
   U8652 : OAI22_X1 port map( A1 => n11208, A2 => n218, B1 => n4921, B2 => n140
                           , ZN => n7889);
   U8653 : AOI22_X1 port map( A1 => n7866, A2 => n4922, B1 => n7867, B2 => 
                           n4923, ZN => n7887);
   U8654 : AOI22_X1 port map( A1 => n7868, A2 => n4924, B1 => n7869, B2 => 
                           n4925, ZN => n7886);
   U8655 : NAND3_X1 port map( A1 => n7890, A2 => n7891, A3 => n7892, ZN => 
                           n12570);
   U8656 : AOI221_X1 port map( B1 => n7862, B2 => n4929, C1 => n7863, C2 => 
                           MEM_IN(6), A => n7893, ZN => n7892);
   U8657 : OAI22_X1 port map( A1 => n11207, A2 => n218, B1 => n4931, B2 => n140
                           , ZN => n7893);
   U8658 : AOI22_X1 port map( A1 => n7866, A2 => n4932, B1 => n7867, B2 => 
                           n4933, ZN => n7891);
   U8659 : AOI22_X1 port map( A1 => n7868, A2 => n4934, B1 => n7869, B2 => 
                           n4935, ZN => n7890);
   U8660 : NAND3_X1 port map( A1 => n7894, A2 => n7895, A3 => n7896, ZN => 
                           n12569);
   U8661 : AOI221_X1 port map( B1 => n7862, B2 => n4939, C1 => n7863, C2 => 
                           MEM_IN(7), A => n7897, ZN => n7896);
   U8662 : OAI22_X1 port map( A1 => n11206, A2 => n218, B1 => n4941, B2 => n140
                           , ZN => n7897);
   U8663 : AOI22_X1 port map( A1 => n7866, A2 => n4942, B1 => n7867, B2 => 
                           n4943, ZN => n7895);
   U8664 : AOI22_X1 port map( A1 => n7868, A2 => n4944, B1 => n7869, B2 => 
                           n4945, ZN => n7894);
   U8665 : NAND3_X1 port map( A1 => n7898, A2 => n7899, A3 => n7900, ZN => 
                           n12568);
   U8666 : AOI221_X1 port map( B1 => n7862, B2 => n4949, C1 => n7863, C2 => 
                           MEM_IN(8), A => n7901, ZN => n7900);
   U8667 : OAI22_X1 port map( A1 => n11205, A2 => n218, B1 => n4951, B2 => n140
                           , ZN => n7901);
   U8668 : AOI22_X1 port map( A1 => n7866, A2 => n4952, B1 => n7867, B2 => 
                           n4953, ZN => n7899);
   U8669 : AOI22_X1 port map( A1 => n7868, A2 => n4954, B1 => n7869, B2 => 
                           n4955, ZN => n7898);
   U8670 : NAND3_X1 port map( A1 => n7902, A2 => n7903, A3 => n7904, ZN => 
                           n12567);
   U8671 : AOI221_X1 port map( B1 => n7862, B2 => n4959, C1 => n7863, C2 => 
                           MEM_IN(9), A => n7905, ZN => n7904);
   U8672 : OAI22_X1 port map( A1 => n11204, A2 => n218, B1 => n4961, B2 => n140
                           , ZN => n7905);
   U8673 : AOI22_X1 port map( A1 => n7866, A2 => n4962, B1 => n7867, B2 => 
                           n4963, ZN => n7903);
   U8674 : AOI22_X1 port map( A1 => n7868, A2 => n4964, B1 => n7869, B2 => 
                           n4965, ZN => n7902);
   U8675 : NAND3_X1 port map( A1 => n7906, A2 => n7907, A3 => n7908, ZN => 
                           n12566);
   U8676 : AOI221_X1 port map( B1 => n7862, B2 => n4969, C1 => n7863, C2 => 
                           MEM_IN(10), A => n7909, ZN => n7908);
   U8677 : OAI22_X1 port map( A1 => n11203, A2 => n218, B1 => n4971, B2 => n140
                           , ZN => n7909);
   U8678 : AOI22_X1 port map( A1 => n7866, A2 => n4972, B1 => n7867, B2 => 
                           n4973, ZN => n7907);
   U8679 : AOI22_X1 port map( A1 => n7868, A2 => n4974, B1 => n7869, B2 => 
                           n4975, ZN => n7906);
   U8680 : NAND3_X1 port map( A1 => n7910, A2 => n7911, A3 => n7912, ZN => 
                           n12565);
   U8681 : AOI221_X1 port map( B1 => n7862, B2 => n4979, C1 => n7863, C2 => 
                           MEM_IN(11), A => n7913, ZN => n7912);
   U8682 : OAI22_X1 port map( A1 => n11202, A2 => n218, B1 => n4981, B2 => n140
                           , ZN => n7913);
   U8683 : AOI22_X1 port map( A1 => n7866, A2 => n4982, B1 => n7867, B2 => 
                           n4983, ZN => n7911);
   U8684 : AOI22_X1 port map( A1 => n7868, A2 => n4984, B1 => n7869, B2 => 
                           n4985, ZN => n7910);
   U8685 : NAND3_X1 port map( A1 => n7914, A2 => n7915, A3 => n7916, ZN => 
                           n12564);
   U8686 : AOI221_X1 port map( B1 => n7862, B2 => n4989, C1 => n7863, C2 => 
                           MEM_IN(12), A => n7917, ZN => n7916);
   U8687 : OAI22_X1 port map( A1 => n11201, A2 => n218, B1 => n4991, B2 => n140
                           , ZN => n7917);
   U8688 : AOI22_X1 port map( A1 => n7866, A2 => n4992, B1 => n7867, B2 => 
                           n4993, ZN => n7915);
   U8689 : AOI22_X1 port map( A1 => n7868, A2 => n4994, B1 => n7869, B2 => 
                           n4995, ZN => n7914);
   U8690 : NAND3_X1 port map( A1 => n7918, A2 => n7919, A3 => n7920, ZN => 
                           n12563);
   U8691 : AOI221_X1 port map( B1 => n7862, B2 => n4999, C1 => n7863, C2 => 
                           MEM_IN(13), A => n7921, ZN => n7920);
   U8692 : OAI22_X1 port map( A1 => n11200, A2 => n218, B1 => n5001, B2 => n140
                           , ZN => n7921);
   U8693 : AOI22_X1 port map( A1 => n7866, A2 => n5002, B1 => n7867, B2 => 
                           n5003, ZN => n7919);
   U8694 : AOI22_X1 port map( A1 => n7868, A2 => n5004, B1 => n7869, B2 => 
                           n5005, ZN => n7918);
   U8695 : NAND3_X1 port map( A1 => n7922, A2 => n7923, A3 => n7924, ZN => 
                           n12562);
   U8696 : AOI221_X1 port map( B1 => n7862, B2 => n5009, C1 => n7863, C2 => 
                           MEM_IN(14), A => n7925, ZN => n7924);
   U8697 : OAI22_X1 port map( A1 => n11199, A2 => n218, B1 => n5011, B2 => n140
                           , ZN => n7925);
   U8698 : AOI22_X1 port map( A1 => n7866, A2 => n5012, B1 => n7867, B2 => 
                           n5013, ZN => n7923);
   U8699 : AOI22_X1 port map( A1 => n7868, A2 => n5014, B1 => n7869, B2 => 
                           n5015, ZN => n7922);
   U8700 : NAND3_X1 port map( A1 => n7926, A2 => n7927, A3 => n7928, ZN => 
                           n12561);
   U8701 : AOI221_X1 port map( B1 => n7862, B2 => n5019, C1 => n7863, C2 => 
                           MEM_IN(15), A => n7929, ZN => n7928);
   U8702 : OAI22_X1 port map( A1 => n11198, A2 => n218, B1 => n5021, B2 => n140
                           , ZN => n7929);
   U8703 : AOI22_X1 port map( A1 => n7866, A2 => n5022, B1 => n7867, B2 => 
                           n5023, ZN => n7927);
   U8704 : AOI22_X1 port map( A1 => n7868, A2 => n5024, B1 => n7869, B2 => 
                           n5025, ZN => n7926);
   U8705 : NAND3_X1 port map( A1 => n7930, A2 => n7931, A3 => n7932, ZN => 
                           n12560);
   U8706 : AOI221_X1 port map( B1 => n7862, B2 => n5029, C1 => n7863, C2 => 
                           MEM_IN(16), A => n7933, ZN => n7932);
   U8707 : OAI22_X1 port map( A1 => n11197, A2 => n218, B1 => n5031, B2 => n140
                           , ZN => n7933);
   U8708 : AOI22_X1 port map( A1 => n7866, A2 => n5032, B1 => n7867, B2 => 
                           n5033, ZN => n7931);
   U8709 : AOI22_X1 port map( A1 => n7868, A2 => n5034, B1 => n7869, B2 => 
                           n5035, ZN => n7930);
   U8710 : NAND3_X1 port map( A1 => n7934, A2 => n7935, A3 => n7936, ZN => 
                           n12559);
   U8711 : AOI221_X1 port map( B1 => n7862, B2 => n5039, C1 => n7863, C2 => 
                           MEM_IN(17), A => n7937, ZN => n7936);
   U8712 : OAI22_X1 port map( A1 => n11196, A2 => n218, B1 => n5041, B2 => n140
                           , ZN => n7937);
   U8713 : AOI22_X1 port map( A1 => n7866, A2 => n5042, B1 => n7867, B2 => 
                           n5043, ZN => n7935);
   U8714 : AOI22_X1 port map( A1 => n7868, A2 => n5044, B1 => n7869, B2 => 
                           n5045, ZN => n7934);
   U8715 : NAND3_X1 port map( A1 => n7938, A2 => n7939, A3 => n7940, ZN => 
                           n12558);
   U8716 : AOI221_X1 port map( B1 => n7862, B2 => n5049, C1 => n7863, C2 => 
                           MEM_IN(18), A => n7941, ZN => n7940);
   U8717 : OAI22_X1 port map( A1 => n11195, A2 => n218, B1 => n5051, B2 => n140
                           , ZN => n7941);
   U8718 : AOI22_X1 port map( A1 => n7866, A2 => n5052, B1 => n7867, B2 => 
                           n5053, ZN => n7939);
   U8719 : AOI22_X1 port map( A1 => n7868, A2 => n5054, B1 => n7869, B2 => 
                           n5055, ZN => n7938);
   U8720 : NAND3_X1 port map( A1 => n7942, A2 => n7943, A3 => n7944, ZN => 
                           n12557);
   U8721 : AOI221_X1 port map( B1 => n7862, B2 => n5059, C1 => n7863, C2 => 
                           MEM_IN(19), A => n7945, ZN => n7944);
   U8722 : OAI22_X1 port map( A1 => n11194, A2 => n218, B1 => n5061, B2 => n140
                           , ZN => n7945);
   U8723 : AOI22_X1 port map( A1 => n7866, A2 => n5062, B1 => n7867, B2 => 
                           n5063, ZN => n7943);
   U8724 : AOI22_X1 port map( A1 => n7868, A2 => n5064, B1 => n7869, B2 => 
                           n5065, ZN => n7942);
   U8725 : NAND3_X1 port map( A1 => n7946, A2 => n7947, A3 => n7948, ZN => 
                           n12556);
   U8726 : AOI221_X1 port map( B1 => n7862, B2 => n5069, C1 => n7863, C2 => 
                           MEM_IN(20), A => n7949, ZN => n7948);
   U8727 : OAI22_X1 port map( A1 => n11193, A2 => n218, B1 => n5071, B2 => n140
                           , ZN => n7949);
   U8728 : AOI22_X1 port map( A1 => n7866, A2 => n5072, B1 => n7867, B2 => 
                           n5073, ZN => n7947);
   U8729 : AOI22_X1 port map( A1 => n7868, A2 => n5074, B1 => n7869, B2 => 
                           n5075, ZN => n7946);
   U8730 : NAND3_X1 port map( A1 => n7950, A2 => n7951, A3 => n7952, ZN => 
                           n12555);
   U8731 : AOI221_X1 port map( B1 => n7862, B2 => n5079, C1 => n7863, C2 => 
                           MEM_IN(21), A => n7953, ZN => n7952);
   U8732 : OAI22_X1 port map( A1 => n11192, A2 => n218, B1 => n5081, B2 => n140
                           , ZN => n7953);
   U8733 : AOI22_X1 port map( A1 => n7866, A2 => n5082, B1 => n7867, B2 => 
                           n5083, ZN => n7951);
   U8734 : AOI22_X1 port map( A1 => n7868, A2 => n5084, B1 => n7869, B2 => 
                           n5085, ZN => n7950);
   U8735 : NAND3_X1 port map( A1 => n7954, A2 => n7955, A3 => n7956, ZN => 
                           n12554);
   U8736 : AOI221_X1 port map( B1 => n7862, B2 => n5089, C1 => n7863, C2 => 
                           MEM_IN(22), A => n7957, ZN => n7956);
   U8737 : OAI22_X1 port map( A1 => n11191, A2 => n218, B1 => n5091, B2 => n140
                           , ZN => n7957);
   U8738 : AOI22_X1 port map( A1 => n7866, A2 => n5092, B1 => n7867, B2 => 
                           n5093, ZN => n7955);
   U8739 : AOI22_X1 port map( A1 => n7868, A2 => n5094, B1 => n7869, B2 => 
                           n5095, ZN => n7954);
   U8740 : NAND3_X1 port map( A1 => n7958, A2 => n7959, A3 => n7960, ZN => 
                           n12553);
   U8741 : AOI221_X1 port map( B1 => n7862, B2 => n5099, C1 => n7863, C2 => 
                           MEM_IN(23), A => n7961, ZN => n7960);
   U8742 : OAI22_X1 port map( A1 => n11190, A2 => n218, B1 => n5101, B2 => n140
                           , ZN => n7961);
   U8743 : AOI22_X1 port map( A1 => n7866, A2 => n5102, B1 => n7867, B2 => 
                           n5103, ZN => n7959);
   U8744 : AOI22_X1 port map( A1 => n7868, A2 => n5104, B1 => n7869, B2 => 
                           n5105, ZN => n7958);
   U8745 : NAND3_X1 port map( A1 => n7962, A2 => n7963, A3 => n7964, ZN => 
                           n12552);
   U8746 : AOI221_X1 port map( B1 => n7862, B2 => n5109, C1 => n7863, C2 => 
                           MEM_IN(24), A => n7965, ZN => n7964);
   U8747 : OAI22_X1 port map( A1 => n11189, A2 => n218, B1 => n5111, B2 => n140
                           , ZN => n7965);
   U8748 : AOI22_X1 port map( A1 => n7866, A2 => n5112, B1 => n7867, B2 => 
                           n5113, ZN => n7963);
   U8749 : AOI22_X1 port map( A1 => n7868, A2 => n5114, B1 => n7869, B2 => 
                           n5115, ZN => n7962);
   U8750 : NAND3_X1 port map( A1 => n7966, A2 => n7967, A3 => n7968, ZN => 
                           n12551);
   U8751 : AOI221_X1 port map( B1 => n7862, B2 => n5119, C1 => n7863, C2 => 
                           MEM_IN(25), A => n7969, ZN => n7968);
   U8752 : OAI22_X1 port map( A1 => n11188, A2 => n218, B1 => n5121, B2 => n140
                           , ZN => n7969);
   U8753 : AOI22_X1 port map( A1 => n7866, A2 => n5122, B1 => n7867, B2 => 
                           n5123, ZN => n7967);
   U8754 : AOI22_X1 port map( A1 => n7868, A2 => n5124, B1 => n7869, B2 => 
                           n5125, ZN => n7966);
   U8755 : NAND3_X1 port map( A1 => n7970, A2 => n7971, A3 => n7972, ZN => 
                           n12550);
   U8756 : AOI221_X1 port map( B1 => n7862, B2 => n5129, C1 => n7863, C2 => 
                           MEM_IN(26), A => n7973, ZN => n7972);
   U8757 : OAI22_X1 port map( A1 => n11187, A2 => n218, B1 => n5131, B2 => n140
                           , ZN => n7973);
   U8758 : AOI22_X1 port map( A1 => n7866, A2 => n5132, B1 => n7867, B2 => 
                           n5133, ZN => n7971);
   U8759 : AOI22_X1 port map( A1 => n7868, A2 => n5134, B1 => n7869, B2 => 
                           n5135, ZN => n7970);
   U8760 : NAND3_X1 port map( A1 => n7974, A2 => n7975, A3 => n7976, ZN => 
                           n12549);
   U8761 : AOI221_X1 port map( B1 => n7862, B2 => n5139, C1 => n7863, C2 => 
                           MEM_IN(27), A => n7977, ZN => n7976);
   U8762 : OAI22_X1 port map( A1 => n11186, A2 => n218, B1 => n5141, B2 => n140
                           , ZN => n7977);
   U8763 : AOI22_X1 port map( A1 => n7866, A2 => n5142, B1 => n7867, B2 => 
                           n5143, ZN => n7975);
   U8764 : AOI22_X1 port map( A1 => n7868, A2 => n5144, B1 => n7869, B2 => 
                           n5145, ZN => n7974);
   U8765 : NAND3_X1 port map( A1 => n7978, A2 => n7979, A3 => n7980, ZN => 
                           n12548);
   U8766 : AOI221_X1 port map( B1 => n7862, B2 => n5149, C1 => n7863, C2 => 
                           MEM_IN(28), A => n7981, ZN => n7980);
   U8767 : OAI22_X1 port map( A1 => n11185, A2 => n218, B1 => n5151, B2 => n140
                           , ZN => n7981);
   U8768 : AOI22_X1 port map( A1 => n7866, A2 => n5152, B1 => n7867, B2 => 
                           n5153, ZN => n7979);
   U8769 : AOI22_X1 port map( A1 => n7868, A2 => n5154, B1 => n7869, B2 => 
                           n5155, ZN => n7978);
   U8770 : NAND3_X1 port map( A1 => n7982, A2 => n7983, A3 => n7984, ZN => 
                           n12547);
   U8771 : AOI221_X1 port map( B1 => n7862, B2 => n5159, C1 => n7863, C2 => 
                           MEM_IN(29), A => n7985, ZN => n7984);
   U8772 : OAI22_X1 port map( A1 => n11184, A2 => n218, B1 => n5161, B2 => n140
                           , ZN => n7985);
   U8773 : AOI22_X1 port map( A1 => n7866, A2 => n5162, B1 => n7867, B2 => 
                           n5163, ZN => n7983);
   U8774 : AOI22_X1 port map( A1 => n7868, A2 => n5164, B1 => n7869, B2 => 
                           n5165, ZN => n7982);
   U8775 : NAND3_X1 port map( A1 => n7986, A2 => n7987, A3 => n7988, ZN => 
                           n12546);
   U8776 : AOI221_X1 port map( B1 => n7862, B2 => n5169, C1 => n7863, C2 => 
                           MEM_IN(30), A => n7989, ZN => n7988);
   U8777 : OAI22_X1 port map( A1 => n11183, A2 => n218, B1 => n5171, B2 => n140
                           , ZN => n7989);
   U8778 : AOI22_X1 port map( A1 => n7866, A2 => n5172, B1 => n7867, B2 => 
                           n5173, ZN => n7987);
   U8779 : AOI22_X1 port map( A1 => n7868, A2 => n5174, B1 => n7869, B2 => 
                           n5175, ZN => n7986);
   U8780 : NAND3_X1 port map( A1 => n7990, A2 => n7991, A3 => n7992, ZN => 
                           n12545);
   U8781 : AOI221_X1 port map( B1 => n7862, B2 => n5179, C1 => n7863, C2 => 
                           MEM_IN(31), A => n7993, ZN => n7992);
   U8782 : OAI22_X1 port map( A1 => n11182, A2 => n218, B1 => n5181, B2 => n140
                           , ZN => n7993);
   U8783 : AOI22_X1 port map( A1 => n7866, A2 => n5191, B1 => n7867, B2 => 
                           n5192, ZN => n7991);
   U8784 : AOI22_X1 port map( A1 => n7868, A2 => n5195, B1 => n7869, B2 => 
                           n5196, ZN => n7990);
   U8785 : OAI22_X1 port map( A1 => n7995, A2 => n7999, B1 => n208, B2 => n217,
                           ZN => n7997);
   U8786 : INV_X1 port map( A => n7994, ZN => n7999);
   U8787 : NOR3_X1 port map( A1 => n4841, A2 => n217, A3 => n6972, ZN => n7994)
                           ;
   U8788 : OAI22_X1 port map( A1 => n4786, A2 => n8000, B1 => n8001, B2 => 
                           n5204, ZN => n7865);
   U8789 : NOR2_X1 port map( A1 => n6972, A2 => n7995, ZN => n8001);
   U8790 : NAND2_X1 port map( A1 => n8002, A2 => n7557, ZN => n6972);
   U8791 : INV_X1 port map( A => n8003, ZN => n7557);
   U8792 : AOI211_X1 port map( C1 => n7705, C2 => n5522, A => n8004, B => RESET
                           , ZN => n8000);
   U8793 : INV_X1 port map( A => n7996, ZN => n8004);
   U8794 : AOI21_X1 port map( B1 => n8003, B2 => n5206, A => n7998, ZN => n7996
                           );
   U8795 : NAND2_X1 port map( A1 => n7410, A2 => n7413, ZN => n8003);
   U8796 : AND2_X1 port map( A1 => n7266, A2 => n7120, ZN => n7410);
   U8797 : NAND2_X1 port map( A1 => n8005, A2 => n8006, ZN => n7995);
   U8798 : NOR2_X1 port map( A1 => n7120, A2 => n4787, ZN => n7554);
   U8799 : NAND2_X1 port map( A1 => n7708, A2 => n5526, ZN => n7120);
   U8800 : NAND3_X1 port map( A1 => n8007, A2 => n8008, A3 => n8009, ZN => 
                           n12544);
   U8801 : AOI221_X1 port map( B1 => n8010, B2 => n4863, C1 => n188, C2 => 
                           MEM_IN(0), A => n8011, ZN => n8009);
   U8802 : OAI22_X1 port map( A1 => n11181, A2 => n265, B1 => n4867, B2 => n141
                           , ZN => n8011);
   U8803 : AOI22_X1 port map( A1 => n200, A2 => n4869, B1 => n8013, B2 => n4871
                           , ZN => n8008);
   U8804 : AOI22_X1 port map( A1 => n242, A2 => n4873, B1 => n8014, B2 => n4875
                           , ZN => n8007);
   U8805 : NAND3_X1 port map( A1 => n8015, A2 => n8016, A3 => n8017, ZN => 
                           n12543);
   U8806 : AOI221_X1 port map( B1 => n8010, B2 => n4879, C1 => n188, C2 => 
                           MEM_IN(1), A => n8018, ZN => n8017);
   U8807 : OAI22_X1 port map( A1 => n11180, A2 => n265, B1 => n4881, B2 => n141
                           , ZN => n8018);
   U8808 : AOI22_X1 port map( A1 => n200, A2 => n4882, B1 => n8013, B2 => n4883
                           , ZN => n8016);
   U8809 : AOI22_X1 port map( A1 => n242, A2 => n4884, B1 => n8014, B2 => n4885
                           , ZN => n8015);
   U8810 : NAND3_X1 port map( A1 => n8019, A2 => n8020, A3 => n8021, ZN => 
                           n12542);
   U8811 : AOI221_X1 port map( B1 => n8010, B2 => n4889, C1 => n188, C2 => 
                           MEM_IN(2), A => n8022, ZN => n8021);
   U8812 : OAI22_X1 port map( A1 => n11179, A2 => n265, B1 => n4891, B2 => n141
                           , ZN => n8022);
   U8813 : AOI22_X1 port map( A1 => n200, A2 => n4892, B1 => n8013, B2 => n4893
                           , ZN => n8020);
   U8814 : AOI22_X1 port map( A1 => n242, A2 => n4894, B1 => n8014, B2 => n4895
                           , ZN => n8019);
   U8815 : NAND3_X1 port map( A1 => n8023, A2 => n8024, A3 => n8025, ZN => 
                           n12541);
   U8816 : AOI221_X1 port map( B1 => n8010, B2 => n4899, C1 => n188, C2 => 
                           MEM_IN(3), A => n8026, ZN => n8025);
   U8817 : OAI22_X1 port map( A1 => n11178, A2 => n265, B1 => n4901, B2 => n141
                           , ZN => n8026);
   U8818 : AOI22_X1 port map( A1 => n200, A2 => n4902, B1 => n8013, B2 => n4903
                           , ZN => n8024);
   U8819 : AOI22_X1 port map( A1 => n242, A2 => n4904, B1 => n8014, B2 => n4905
                           , ZN => n8023);
   U8820 : NAND3_X1 port map( A1 => n8027, A2 => n8028, A3 => n8029, ZN => 
                           n12540);
   U8821 : AOI221_X1 port map( B1 => n8010, B2 => n4909, C1 => n188, C2 => 
                           MEM_IN(4), A => n8030, ZN => n8029);
   U8822 : OAI22_X1 port map( A1 => n11177, A2 => n265, B1 => n4911, B2 => n141
                           , ZN => n8030);
   U8823 : AOI22_X1 port map( A1 => n200, A2 => n4912, B1 => n8013, B2 => n4913
                           , ZN => n8028);
   U8824 : AOI22_X1 port map( A1 => n242, A2 => n4914, B1 => n8014, B2 => n4915
                           , ZN => n8027);
   U8825 : NAND3_X1 port map( A1 => n8031, A2 => n8032, A3 => n8033, ZN => 
                           n12539);
   U8826 : AOI221_X1 port map( B1 => n8010, B2 => n4919, C1 => n188, C2 => 
                           MEM_IN(5), A => n8034, ZN => n8033);
   U8827 : OAI22_X1 port map( A1 => n11176, A2 => n265, B1 => n4921, B2 => n141
                           , ZN => n8034);
   U8828 : AOI22_X1 port map( A1 => n200, A2 => n4922, B1 => n8013, B2 => n4923
                           , ZN => n8032);
   U8829 : AOI22_X1 port map( A1 => n242, A2 => n4924, B1 => n8014, B2 => n4925
                           , ZN => n8031);
   U8830 : NAND3_X1 port map( A1 => n8035, A2 => n8036, A3 => n8037, ZN => 
                           n12538);
   U8831 : AOI221_X1 port map( B1 => n8010, B2 => n4929, C1 => n188, C2 => 
                           MEM_IN(6), A => n8038, ZN => n8037);
   U8832 : OAI22_X1 port map( A1 => n11175, A2 => n265, B1 => n4931, B2 => n141
                           , ZN => n8038);
   U8833 : AOI22_X1 port map( A1 => n200, A2 => n4932, B1 => n8013, B2 => n4933
                           , ZN => n8036);
   U8834 : AOI22_X1 port map( A1 => n242, A2 => n4934, B1 => n8014, B2 => n4935
                           , ZN => n8035);
   U8835 : NAND3_X1 port map( A1 => n8039, A2 => n8040, A3 => n8041, ZN => 
                           n12537);
   U8836 : AOI221_X1 port map( B1 => n8010, B2 => n4939, C1 => n188, C2 => 
                           MEM_IN(7), A => n8042, ZN => n8041);
   U8837 : OAI22_X1 port map( A1 => n11174, A2 => n265, B1 => n4941, B2 => n141
                           , ZN => n8042);
   U8838 : AOI22_X1 port map( A1 => n200, A2 => n4942, B1 => n8013, B2 => n4943
                           , ZN => n8040);
   U8839 : AOI22_X1 port map( A1 => n242, A2 => n4944, B1 => n8014, B2 => n4945
                           , ZN => n8039);
   U8840 : NAND3_X1 port map( A1 => n8043, A2 => n8044, A3 => n8045, ZN => 
                           n12536);
   U8841 : AOI221_X1 port map( B1 => n8010, B2 => n4949, C1 => n188, C2 => 
                           MEM_IN(8), A => n8046, ZN => n8045);
   U8842 : OAI22_X1 port map( A1 => n11173, A2 => n265, B1 => n4951, B2 => n141
                           , ZN => n8046);
   U8843 : AOI22_X1 port map( A1 => n200, A2 => n4952, B1 => n8013, B2 => n4953
                           , ZN => n8044);
   U8844 : AOI22_X1 port map( A1 => n242, A2 => n4954, B1 => n8014, B2 => n4955
                           , ZN => n8043);
   U8845 : NAND3_X1 port map( A1 => n8047, A2 => n8048, A3 => n8049, ZN => 
                           n12535);
   U8846 : AOI221_X1 port map( B1 => n8010, B2 => n4959, C1 => n188, C2 => 
                           MEM_IN(9), A => n8050, ZN => n8049);
   U8847 : OAI22_X1 port map( A1 => n11172, A2 => n265, B1 => n4961, B2 => n141
                           , ZN => n8050);
   U8848 : AOI22_X1 port map( A1 => n200, A2 => n4962, B1 => n8013, B2 => n4963
                           , ZN => n8048);
   U8849 : AOI22_X1 port map( A1 => n242, A2 => n4964, B1 => n8014, B2 => n4965
                           , ZN => n8047);
   U8850 : NAND3_X1 port map( A1 => n8051, A2 => n8052, A3 => n8053, ZN => 
                           n12534);
   U8851 : AOI221_X1 port map( B1 => n8010, B2 => n4969, C1 => n188, C2 => 
                           MEM_IN(10), A => n8054, ZN => n8053);
   U8852 : OAI22_X1 port map( A1 => n11171, A2 => n265, B1 => n4971, B2 => n141
                           , ZN => n8054);
   U8853 : AOI22_X1 port map( A1 => n200, A2 => n4972, B1 => n8013, B2 => n4973
                           , ZN => n8052);
   U8854 : AOI22_X1 port map( A1 => n242, A2 => n4974, B1 => n8014, B2 => n4975
                           , ZN => n8051);
   U8855 : NAND3_X1 port map( A1 => n8055, A2 => n8056, A3 => n8057, ZN => 
                           n12533);
   U8856 : AOI221_X1 port map( B1 => n8010, B2 => n4979, C1 => n188, C2 => 
                           MEM_IN(11), A => n8058, ZN => n8057);
   U8857 : OAI22_X1 port map( A1 => n11170, A2 => n265, B1 => n4981, B2 => n141
                           , ZN => n8058);
   U8858 : AOI22_X1 port map( A1 => n200, A2 => n4982, B1 => n8013, B2 => n4983
                           , ZN => n8056);
   U8859 : AOI22_X1 port map( A1 => n242, A2 => n4984, B1 => n8014, B2 => n4985
                           , ZN => n8055);
   U8860 : NAND3_X1 port map( A1 => n8059, A2 => n8060, A3 => n8061, ZN => 
                           n12532);
   U8861 : AOI221_X1 port map( B1 => n8010, B2 => n4989, C1 => n188, C2 => 
                           MEM_IN(12), A => n8062, ZN => n8061);
   U8862 : OAI22_X1 port map( A1 => n11169, A2 => n265, B1 => n4991, B2 => n141
                           , ZN => n8062);
   U8863 : AOI22_X1 port map( A1 => n200, A2 => n4992, B1 => n8013, B2 => n4993
                           , ZN => n8060);
   U8864 : AOI22_X1 port map( A1 => n242, A2 => n4994, B1 => n8014, B2 => n4995
                           , ZN => n8059);
   U8865 : NAND3_X1 port map( A1 => n8063, A2 => n8064, A3 => n8065, ZN => 
                           n12531);
   U8866 : AOI221_X1 port map( B1 => n8010, B2 => n4999, C1 => n188, C2 => 
                           MEM_IN(13), A => n8066, ZN => n8065);
   U8867 : OAI22_X1 port map( A1 => n11168, A2 => n265, B1 => n5001, B2 => n141
                           , ZN => n8066);
   U8868 : AOI22_X1 port map( A1 => n200, A2 => n5002, B1 => n8013, B2 => n5003
                           , ZN => n8064);
   U8869 : AOI22_X1 port map( A1 => n242, A2 => n5004, B1 => n8014, B2 => n5005
                           , ZN => n8063);
   U8870 : NAND3_X1 port map( A1 => n8067, A2 => n8068, A3 => n8069, ZN => 
                           n12530);
   U8871 : AOI221_X1 port map( B1 => n8010, B2 => n5009, C1 => n188, C2 => 
                           MEM_IN(14), A => n8070, ZN => n8069);
   U8872 : OAI22_X1 port map( A1 => n11167, A2 => n265, B1 => n5011, B2 => n141
                           , ZN => n8070);
   U8873 : AOI22_X1 port map( A1 => n200, A2 => n5012, B1 => n8013, B2 => n5013
                           , ZN => n8068);
   U8874 : AOI22_X1 port map( A1 => n242, A2 => n5014, B1 => n8014, B2 => n5015
                           , ZN => n8067);
   U8875 : NAND3_X1 port map( A1 => n8071, A2 => n8072, A3 => n8073, ZN => 
                           n12529);
   U8876 : AOI221_X1 port map( B1 => n8010, B2 => n5019, C1 => n188, C2 => 
                           MEM_IN(15), A => n8074, ZN => n8073);
   U8877 : OAI22_X1 port map( A1 => n11166, A2 => n265, B1 => n5021, B2 => n141
                           , ZN => n8074);
   U8878 : AOI22_X1 port map( A1 => n200, A2 => n5022, B1 => n8013, B2 => n5023
                           , ZN => n8072);
   U8879 : AOI22_X1 port map( A1 => n242, A2 => n5024, B1 => n8014, B2 => n5025
                           , ZN => n8071);
   U8880 : NAND3_X1 port map( A1 => n8075, A2 => n8076, A3 => n8077, ZN => 
                           n12528);
   U8881 : AOI221_X1 port map( B1 => n8010, B2 => n5029, C1 => n188, C2 => 
                           MEM_IN(16), A => n8078, ZN => n8077);
   U8882 : OAI22_X1 port map( A1 => n11165, A2 => n265, B1 => n5031, B2 => n141
                           , ZN => n8078);
   U8883 : AOI22_X1 port map( A1 => n200, A2 => n5032, B1 => n8013, B2 => n5033
                           , ZN => n8076);
   U8884 : AOI22_X1 port map( A1 => n242, A2 => n5034, B1 => n8014, B2 => n5035
                           , ZN => n8075);
   U8885 : NAND3_X1 port map( A1 => n8079, A2 => n8080, A3 => n8081, ZN => 
                           n12527);
   U8886 : AOI221_X1 port map( B1 => n8010, B2 => n5039, C1 => n188, C2 => 
                           MEM_IN(17), A => n8082, ZN => n8081);
   U8887 : OAI22_X1 port map( A1 => n11164, A2 => n265, B1 => n5041, B2 => n141
                           , ZN => n8082);
   U8888 : AOI22_X1 port map( A1 => n200, A2 => n5042, B1 => n8013, B2 => n5043
                           , ZN => n8080);
   U8889 : AOI22_X1 port map( A1 => n242, A2 => n5044, B1 => n8014, B2 => n5045
                           , ZN => n8079);
   U8890 : NAND3_X1 port map( A1 => n8083, A2 => n8084, A3 => n8085, ZN => 
                           n12526);
   U8891 : AOI221_X1 port map( B1 => n8010, B2 => n5049, C1 => n188, C2 => 
                           MEM_IN(18), A => n8086, ZN => n8085);
   U8892 : OAI22_X1 port map( A1 => n11163, A2 => n265, B1 => n5051, B2 => n141
                           , ZN => n8086);
   U8893 : AOI22_X1 port map( A1 => n200, A2 => n5052, B1 => n8013, B2 => n5053
                           , ZN => n8084);
   U8894 : AOI22_X1 port map( A1 => n242, A2 => n5054, B1 => n8014, B2 => n5055
                           , ZN => n8083);
   U8895 : NAND3_X1 port map( A1 => n8087, A2 => n8088, A3 => n8089, ZN => 
                           n12525);
   U8896 : AOI221_X1 port map( B1 => n8010, B2 => n5059, C1 => n188, C2 => 
                           MEM_IN(19), A => n8090, ZN => n8089);
   U8897 : OAI22_X1 port map( A1 => n11162, A2 => n265, B1 => n5061, B2 => n141
                           , ZN => n8090);
   U8898 : AOI22_X1 port map( A1 => n200, A2 => n5062, B1 => n8013, B2 => n5063
                           , ZN => n8088);
   U8899 : AOI22_X1 port map( A1 => n242, A2 => n5064, B1 => n8014, B2 => n5065
                           , ZN => n8087);
   U8900 : NAND3_X1 port map( A1 => n8091, A2 => n8092, A3 => n8093, ZN => 
                           n12524);
   U8901 : AOI221_X1 port map( B1 => n8010, B2 => n5069, C1 => n188, C2 => 
                           MEM_IN(20), A => n8094, ZN => n8093);
   U8902 : OAI22_X1 port map( A1 => n11161, A2 => n265, B1 => n5071, B2 => n141
                           , ZN => n8094);
   U8903 : AOI22_X1 port map( A1 => n200, A2 => n5072, B1 => n8013, B2 => n5073
                           , ZN => n8092);
   U8904 : AOI22_X1 port map( A1 => n242, A2 => n5074, B1 => n8014, B2 => n5075
                           , ZN => n8091);
   U8905 : NAND3_X1 port map( A1 => n8095, A2 => n8096, A3 => n8097, ZN => 
                           n12523);
   U8906 : AOI221_X1 port map( B1 => n8010, B2 => n5079, C1 => n188, C2 => 
                           MEM_IN(21), A => n8098, ZN => n8097);
   U8907 : OAI22_X1 port map( A1 => n11160, A2 => n265, B1 => n5081, B2 => n141
                           , ZN => n8098);
   U8908 : AOI22_X1 port map( A1 => n200, A2 => n5082, B1 => n8013, B2 => n5083
                           , ZN => n8096);
   U8909 : AOI22_X1 port map( A1 => n242, A2 => n5084, B1 => n8014, B2 => n5085
                           , ZN => n8095);
   U8910 : NAND3_X1 port map( A1 => n8099, A2 => n8100, A3 => n8101, ZN => 
                           n12522);
   U8911 : AOI221_X1 port map( B1 => n8010, B2 => n5089, C1 => n188, C2 => 
                           MEM_IN(22), A => n8102, ZN => n8101);
   U8912 : OAI22_X1 port map( A1 => n11159, A2 => n265, B1 => n5091, B2 => n141
                           , ZN => n8102);
   U8913 : AOI22_X1 port map( A1 => n200, A2 => n5092, B1 => n8013, B2 => n5093
                           , ZN => n8100);
   U8914 : AOI22_X1 port map( A1 => n242, A2 => n5094, B1 => n8014, B2 => n5095
                           , ZN => n8099);
   U8915 : NAND3_X1 port map( A1 => n8103, A2 => n8104, A3 => n8105, ZN => 
                           n12521);
   U8916 : AOI221_X1 port map( B1 => n8010, B2 => n5099, C1 => n188, C2 => 
                           MEM_IN(23), A => n8106, ZN => n8105);
   U8917 : OAI22_X1 port map( A1 => n11158, A2 => n265, B1 => n5101, B2 => n141
                           , ZN => n8106);
   U8918 : AOI22_X1 port map( A1 => n200, A2 => n5102, B1 => n8013, B2 => n5103
                           , ZN => n8104);
   U8919 : AOI22_X1 port map( A1 => n242, A2 => n5104, B1 => n8014, B2 => n5105
                           , ZN => n8103);
   U8920 : NAND3_X1 port map( A1 => n8107, A2 => n8108, A3 => n8109, ZN => 
                           n12520);
   U8921 : AOI221_X1 port map( B1 => n8010, B2 => n5109, C1 => n188, C2 => 
                           MEM_IN(24), A => n8110, ZN => n8109);
   U8922 : OAI22_X1 port map( A1 => n11157, A2 => n265, B1 => n5111, B2 => n141
                           , ZN => n8110);
   U8923 : AOI22_X1 port map( A1 => n200, A2 => n5112, B1 => n8013, B2 => n5113
                           , ZN => n8108);
   U8924 : AOI22_X1 port map( A1 => n242, A2 => n5114, B1 => n8014, B2 => n5115
                           , ZN => n8107);
   U8925 : NAND3_X1 port map( A1 => n8111, A2 => n8112, A3 => n8113, ZN => 
                           n12519);
   U8926 : AOI221_X1 port map( B1 => n8010, B2 => n5119, C1 => n188, C2 => 
                           MEM_IN(25), A => n8114, ZN => n8113);
   U8927 : OAI22_X1 port map( A1 => n11156, A2 => n265, B1 => n5121, B2 => n141
                           , ZN => n8114);
   U8928 : AOI22_X1 port map( A1 => n200, A2 => n5122, B1 => n8013, B2 => n5123
                           , ZN => n8112);
   U8929 : AOI22_X1 port map( A1 => n242, A2 => n5124, B1 => n8014, B2 => n5125
                           , ZN => n8111);
   U8930 : NAND3_X1 port map( A1 => n8115, A2 => n8116, A3 => n8117, ZN => 
                           n12518);
   U8931 : AOI221_X1 port map( B1 => n8010, B2 => n5129, C1 => n188, C2 => 
                           MEM_IN(26), A => n8118, ZN => n8117);
   U8932 : OAI22_X1 port map( A1 => n11155, A2 => n265, B1 => n5131, B2 => n141
                           , ZN => n8118);
   U8933 : AOI22_X1 port map( A1 => n200, A2 => n5132, B1 => n8013, B2 => n5133
                           , ZN => n8116);
   U8934 : AOI22_X1 port map( A1 => n242, A2 => n5134, B1 => n8014, B2 => n5135
                           , ZN => n8115);
   U8935 : NAND3_X1 port map( A1 => n8119, A2 => n8120, A3 => n8121, ZN => 
                           n12517);
   U8936 : AOI221_X1 port map( B1 => n8010, B2 => n5139, C1 => n188, C2 => 
                           MEM_IN(27), A => n8122, ZN => n8121);
   U8937 : OAI22_X1 port map( A1 => n11154, A2 => n265, B1 => n5141, B2 => n141
                           , ZN => n8122);
   U8938 : AOI22_X1 port map( A1 => n200, A2 => n5142, B1 => n8013, B2 => n5143
                           , ZN => n8120);
   U8939 : AOI22_X1 port map( A1 => n242, A2 => n5144, B1 => n8014, B2 => n5145
                           , ZN => n8119);
   U8940 : NAND3_X1 port map( A1 => n8123, A2 => n8124, A3 => n8125, ZN => 
                           n12516);
   U8941 : AOI221_X1 port map( B1 => n8010, B2 => n5149, C1 => n188, C2 => 
                           MEM_IN(28), A => n8126, ZN => n8125);
   U8942 : OAI22_X1 port map( A1 => n11153, A2 => n265, B1 => n5151, B2 => n141
                           , ZN => n8126);
   U8943 : AOI22_X1 port map( A1 => n200, A2 => n5152, B1 => n8013, B2 => n5153
                           , ZN => n8124);
   U8944 : AOI22_X1 port map( A1 => n242, A2 => n5154, B1 => n8014, B2 => n5155
                           , ZN => n8123);
   U8945 : NAND3_X1 port map( A1 => n8127, A2 => n8128, A3 => n8129, ZN => 
                           n12515);
   U8946 : AOI221_X1 port map( B1 => n8010, B2 => n5159, C1 => n188, C2 => 
                           MEM_IN(29), A => n8130, ZN => n8129);
   U8947 : OAI22_X1 port map( A1 => n11152, A2 => n265, B1 => n5161, B2 => n141
                           , ZN => n8130);
   U8948 : AOI22_X1 port map( A1 => n200, A2 => n5162, B1 => n8013, B2 => n5163
                           , ZN => n8128);
   U8949 : AOI22_X1 port map( A1 => n242, A2 => n5164, B1 => n8014, B2 => n5165
                           , ZN => n8127);
   U8950 : NAND3_X1 port map( A1 => n8131, A2 => n8132, A3 => n8133, ZN => 
                           n12514);
   U8951 : AOI221_X1 port map( B1 => n8010, B2 => n5169, C1 => n188, C2 => 
                           MEM_IN(30), A => n8134, ZN => n8133);
   U8952 : OAI22_X1 port map( A1 => n11151, A2 => n265, B1 => n5171, B2 => n141
                           , ZN => n8134);
   U8953 : AOI22_X1 port map( A1 => n200, A2 => n5172, B1 => n8013, B2 => n5173
                           , ZN => n8132);
   U8954 : AOI22_X1 port map( A1 => n242, A2 => n5174, B1 => n8014, B2 => n5175
                           , ZN => n8131);
   U8955 : NAND3_X1 port map( A1 => n8135, A2 => n8136, A3 => n8137, ZN => 
                           n12513);
   U8956 : AOI221_X1 port map( B1 => n8010, B2 => n5179, C1 => n188, C2 => 
                           MEM_IN(31), A => n8138, ZN => n8137);
   U8957 : OAI22_X1 port map( A1 => n11150, A2 => n265, B1 => n5181, B2 => n141
                           , ZN => n8138);
   U8958 : AOI22_X1 port map( A1 => n200, A2 => n5191, B1 => n8013, B2 => n5192
                           , ZN => n8136);
   U8959 : AOI22_X1 port map( A1 => n242, A2 => n5195, B1 => n8014, B2 => n5196
                           , ZN => n8135);
   U8960 : INV_X1 port map( A => n8145, ZN => n8143);
   U8961 : AOI22_X1 port map( A1 => n8141, A2 => n8148, B1 => n4841, B2 => n265
                           , ZN => n8145);
   U8962 : INV_X1 port map( A => n8140, ZN => n8148);
   U8963 : NAND3_X1 port map( A1 => n208, A2 => n265, A3 => n7119, ZN => n8140)
                           ;
   U8964 : INV_X1 port map( A => n8139, ZN => n7119);
   U8965 : OAI22_X1 port map( A1 => n8149, A2 => n4786, B1 => n8150, B2 => 
                           n5204, ZN => n8012);
   U8966 : NOR2_X1 port map( A1 => n8139, A2 => n8151, ZN => n8150);
   U8967 : NAND4_X1 port map( A1 => n8002, A2 => n8006, A3 => n7413, A4 => 
                           n7266, ZN => n8139);
   U8968 : NOR4_X1 port map( A1 => n8152, A2 => n7998, A3 => RESET, A4 => n8153
                           , ZN => n8149);
   U8969 : OAI211_X1 port map( C1 => n5771, C2 => n7856, A => n7698, B => n7847
                           , ZN => n8152);
   U8970 : INV_X1 port map( A => n7849, ZN => n7698);
   U8971 : NOR2_X1 port map( A1 => n7266, A2 => n4787, ZN => n7849);
   U8972 : INV_X1 port map( A => n8151, ZN => n8141);
   U8973 : NAND2_X1 port map( A1 => n8154, A2 => n8155, ZN => n8151);
   U8974 : NAND2_X1 port map( A1 => n7708, A2 => n5775, ZN => n7266);
   U8975 : NAND3_X1 port map( A1 => n8156, A2 => n8157, A3 => n8158, ZN => 
                           n12512);
   U8976 : AOI221_X1 port map( B1 => n8159, B2 => n4863, C1 => n189, C2 => 
                           MEM_IN(0), A => n8160, ZN => n8158);
   U8977 : OAI22_X1 port map( A1 => n11149, A2 => n287, B1 => n4867, B2 => n138
                           , ZN => n8160);
   U8978 : AOI22_X1 port map( A1 => n8162, A2 => n4869, B1 => n8163, B2 => 
                           n4871, ZN => n8157);
   U8979 : AOI22_X1 port map( A1 => n8164, A2 => n4873, B1 => n8165, B2 => 
                           n4875, ZN => n8156);
   U8980 : NAND3_X1 port map( A1 => n8166, A2 => n8167, A3 => n8168, ZN => 
                           n12511);
   U8981 : AOI221_X1 port map( B1 => n8159, B2 => n4879, C1 => n189, C2 => 
                           MEM_IN(1), A => n8169, ZN => n8168);
   U8982 : OAI22_X1 port map( A1 => n11148, A2 => n287, B1 => n4881, B2 => n138
                           , ZN => n8169);
   U8983 : AOI22_X1 port map( A1 => n8162, A2 => n4882, B1 => n8163, B2 => 
                           n4883, ZN => n8167);
   U8984 : AOI22_X1 port map( A1 => n8164, A2 => n4884, B1 => n8165, B2 => 
                           n4885, ZN => n8166);
   U8985 : NAND3_X1 port map( A1 => n8170, A2 => n8171, A3 => n8172, ZN => 
                           n12510);
   U8986 : AOI221_X1 port map( B1 => n8159, B2 => n4889, C1 => n189, C2 => 
                           MEM_IN(2), A => n8173, ZN => n8172);
   U8987 : OAI22_X1 port map( A1 => n11147, A2 => n287, B1 => n4891, B2 => n138
                           , ZN => n8173);
   U8988 : AOI22_X1 port map( A1 => n8162, A2 => n4892, B1 => n8163, B2 => 
                           n4893, ZN => n8171);
   U8989 : AOI22_X1 port map( A1 => n8164, A2 => n4894, B1 => n8165, B2 => 
                           n4895, ZN => n8170);
   U8990 : NAND3_X1 port map( A1 => n8174, A2 => n8175, A3 => n8176, ZN => 
                           n12509);
   U8991 : AOI221_X1 port map( B1 => n8159, B2 => n4899, C1 => n189, C2 => 
                           MEM_IN(3), A => n8177, ZN => n8176);
   U8992 : OAI22_X1 port map( A1 => n11146, A2 => n287, B1 => n4901, B2 => n138
                           , ZN => n8177);
   U8993 : AOI22_X1 port map( A1 => n8162, A2 => n4902, B1 => n8163, B2 => 
                           n4903, ZN => n8175);
   U8994 : AOI22_X1 port map( A1 => n8164, A2 => n4904, B1 => n8165, B2 => 
                           n4905, ZN => n8174);
   U8995 : NAND3_X1 port map( A1 => n8178, A2 => n8179, A3 => n8180, ZN => 
                           n12508);
   U8996 : AOI221_X1 port map( B1 => n8159, B2 => n4909, C1 => n189, C2 => 
                           MEM_IN(4), A => n8181, ZN => n8180);
   U8997 : OAI22_X1 port map( A1 => n11145, A2 => n287, B1 => n4911, B2 => n138
                           , ZN => n8181);
   U8998 : AOI22_X1 port map( A1 => n8162, A2 => n4912, B1 => n8163, B2 => 
                           n4913, ZN => n8179);
   U8999 : AOI22_X1 port map( A1 => n8164, A2 => n4914, B1 => n8165, B2 => 
                           n4915, ZN => n8178);
   U9000 : NAND3_X1 port map( A1 => n8182, A2 => n8183, A3 => n8184, ZN => 
                           n12507);
   U9001 : AOI221_X1 port map( B1 => n8159, B2 => n4919, C1 => n189, C2 => 
                           MEM_IN(5), A => n8185, ZN => n8184);
   U9002 : OAI22_X1 port map( A1 => n11144, A2 => n287, B1 => n4921, B2 => n138
                           , ZN => n8185);
   U9003 : AOI22_X1 port map( A1 => n8162, A2 => n4922, B1 => n8163, B2 => 
                           n4923, ZN => n8183);
   U9004 : AOI22_X1 port map( A1 => n8164, A2 => n4924, B1 => n8165, B2 => 
                           n4925, ZN => n8182);
   U9005 : NAND3_X1 port map( A1 => n8186, A2 => n8187, A3 => n8188, ZN => 
                           n12506);
   U9006 : AOI221_X1 port map( B1 => n8159, B2 => n4929, C1 => n189, C2 => 
                           MEM_IN(6), A => n8189, ZN => n8188);
   U9007 : OAI22_X1 port map( A1 => n11143, A2 => n287, B1 => n4931, B2 => n138
                           , ZN => n8189);
   U9008 : AOI22_X1 port map( A1 => n8162, A2 => n4932, B1 => n8163, B2 => 
                           n4933, ZN => n8187);
   U9009 : AOI22_X1 port map( A1 => n8164, A2 => n4934, B1 => n8165, B2 => 
                           n4935, ZN => n8186);
   U9010 : NAND3_X1 port map( A1 => n8190, A2 => n8191, A3 => n8192, ZN => 
                           n12505);
   U9011 : AOI221_X1 port map( B1 => n8159, B2 => n4939, C1 => n189, C2 => 
                           MEM_IN(7), A => n8193, ZN => n8192);
   U9012 : OAI22_X1 port map( A1 => n11142, A2 => n287, B1 => n4941, B2 => n138
                           , ZN => n8193);
   U9013 : AOI22_X1 port map( A1 => n8162, A2 => n4942, B1 => n8163, B2 => 
                           n4943, ZN => n8191);
   U9014 : AOI22_X1 port map( A1 => n8164, A2 => n4944, B1 => n8165, B2 => 
                           n4945, ZN => n8190);
   U9015 : NAND3_X1 port map( A1 => n8194, A2 => n8195, A3 => n8196, ZN => 
                           n12504);
   U9016 : AOI221_X1 port map( B1 => n8159, B2 => n4949, C1 => n189, C2 => 
                           MEM_IN(8), A => n8197, ZN => n8196);
   U9017 : OAI22_X1 port map( A1 => n11141, A2 => n287, B1 => n4951, B2 => n138
                           , ZN => n8197);
   U9018 : AOI22_X1 port map( A1 => n8162, A2 => n4952, B1 => n8163, B2 => 
                           n4953, ZN => n8195);
   U9019 : AOI22_X1 port map( A1 => n8164, A2 => n4954, B1 => n8165, B2 => 
                           n4955, ZN => n8194);
   U9020 : NAND3_X1 port map( A1 => n8198, A2 => n8199, A3 => n8200, ZN => 
                           n12503);
   U9021 : AOI221_X1 port map( B1 => n8159, B2 => n4959, C1 => n189, C2 => 
                           MEM_IN(9), A => n8201, ZN => n8200);
   U9022 : OAI22_X1 port map( A1 => n11140, A2 => n287, B1 => n4961, B2 => n138
                           , ZN => n8201);
   U9023 : AOI22_X1 port map( A1 => n8162, A2 => n4962, B1 => n8163, B2 => 
                           n4963, ZN => n8199);
   U9024 : AOI22_X1 port map( A1 => n8164, A2 => n4964, B1 => n8165, B2 => 
                           n4965, ZN => n8198);
   U9025 : NAND3_X1 port map( A1 => n8202, A2 => n8203, A3 => n8204, ZN => 
                           n12502);
   U9026 : AOI221_X1 port map( B1 => n8159, B2 => n4969, C1 => n189, C2 => 
                           MEM_IN(10), A => n8205, ZN => n8204);
   U9027 : OAI22_X1 port map( A1 => n11139, A2 => n287, B1 => n4971, B2 => n138
                           , ZN => n8205);
   U9028 : AOI22_X1 port map( A1 => n8162, A2 => n4972, B1 => n8163, B2 => 
                           n4973, ZN => n8203);
   U9029 : AOI22_X1 port map( A1 => n8164, A2 => n4974, B1 => n8165, B2 => 
                           n4975, ZN => n8202);
   U9030 : NAND3_X1 port map( A1 => n8206, A2 => n8207, A3 => n8208, ZN => 
                           n12501);
   U9031 : AOI221_X1 port map( B1 => n8159, B2 => n4979, C1 => n189, C2 => 
                           MEM_IN(11), A => n8209, ZN => n8208);
   U9032 : OAI22_X1 port map( A1 => n11138, A2 => n287, B1 => n4981, B2 => n138
                           , ZN => n8209);
   U9033 : AOI22_X1 port map( A1 => n8162, A2 => n4982, B1 => n8163, B2 => 
                           n4983, ZN => n8207);
   U9034 : AOI22_X1 port map( A1 => n8164, A2 => n4984, B1 => n8165, B2 => 
                           n4985, ZN => n8206);
   U9035 : NAND3_X1 port map( A1 => n8210, A2 => n8211, A3 => n8212, ZN => 
                           n12500);
   U9036 : AOI221_X1 port map( B1 => n8159, B2 => n4989, C1 => n189, C2 => 
                           MEM_IN(12), A => n8213, ZN => n8212);
   U9037 : OAI22_X1 port map( A1 => n11137, A2 => n287, B1 => n4991, B2 => n138
                           , ZN => n8213);
   U9038 : AOI22_X1 port map( A1 => n8162, A2 => n4992, B1 => n8163, B2 => 
                           n4993, ZN => n8211);
   U9039 : AOI22_X1 port map( A1 => n8164, A2 => n4994, B1 => n8165, B2 => 
                           n4995, ZN => n8210);
   U9040 : NAND3_X1 port map( A1 => n8214, A2 => n8215, A3 => n8216, ZN => 
                           n12499);
   U9041 : AOI221_X1 port map( B1 => n8159, B2 => n4999, C1 => n189, C2 => 
                           MEM_IN(13), A => n8217, ZN => n8216);
   U9042 : OAI22_X1 port map( A1 => n11136, A2 => n287, B1 => n5001, B2 => n138
                           , ZN => n8217);
   U9043 : AOI22_X1 port map( A1 => n8162, A2 => n5002, B1 => n8163, B2 => 
                           n5003, ZN => n8215);
   U9044 : AOI22_X1 port map( A1 => n8164, A2 => n5004, B1 => n8165, B2 => 
                           n5005, ZN => n8214);
   U9045 : NAND3_X1 port map( A1 => n8218, A2 => n8219, A3 => n8220, ZN => 
                           n12498);
   U9046 : AOI221_X1 port map( B1 => n8159, B2 => n5009, C1 => n189, C2 => 
                           MEM_IN(14), A => n8221, ZN => n8220);
   U9047 : OAI22_X1 port map( A1 => n11135, A2 => n287, B1 => n5011, B2 => n138
                           , ZN => n8221);
   U9048 : AOI22_X1 port map( A1 => n8162, A2 => n5012, B1 => n8163, B2 => 
                           n5013, ZN => n8219);
   U9049 : AOI22_X1 port map( A1 => n8164, A2 => n5014, B1 => n8165, B2 => 
                           n5015, ZN => n8218);
   U9050 : NAND3_X1 port map( A1 => n8222, A2 => n8223, A3 => n8224, ZN => 
                           n12497);
   U9051 : AOI221_X1 port map( B1 => n8159, B2 => n5019, C1 => n189, C2 => 
                           MEM_IN(15), A => n8225, ZN => n8224);
   U9052 : OAI22_X1 port map( A1 => n11134, A2 => n287, B1 => n5021, B2 => n138
                           , ZN => n8225);
   U9053 : AOI22_X1 port map( A1 => n8162, A2 => n5022, B1 => n8163, B2 => 
                           n5023, ZN => n8223);
   U9054 : AOI22_X1 port map( A1 => n8164, A2 => n5024, B1 => n8165, B2 => 
                           n5025, ZN => n8222);
   U9055 : NAND3_X1 port map( A1 => n8226, A2 => n8227, A3 => n8228, ZN => 
                           n12496);
   U9056 : AOI221_X1 port map( B1 => n8159, B2 => n5029, C1 => n189, C2 => 
                           MEM_IN(16), A => n8229, ZN => n8228);
   U9057 : OAI22_X1 port map( A1 => n11133, A2 => n287, B1 => n5031, B2 => n138
                           , ZN => n8229);
   U9058 : AOI22_X1 port map( A1 => n8162, A2 => n5032, B1 => n8163, B2 => 
                           n5033, ZN => n8227);
   U9059 : AOI22_X1 port map( A1 => n8164, A2 => n5034, B1 => n8165, B2 => 
                           n5035, ZN => n8226);
   U9060 : NAND3_X1 port map( A1 => n8230, A2 => n8231, A3 => n8232, ZN => 
                           n12495);
   U9061 : AOI221_X1 port map( B1 => n8159, B2 => n5039, C1 => n189, C2 => 
                           MEM_IN(17), A => n8233, ZN => n8232);
   U9062 : OAI22_X1 port map( A1 => n11132, A2 => n287, B1 => n5041, B2 => n138
                           , ZN => n8233);
   U9063 : AOI22_X1 port map( A1 => n8162, A2 => n5042, B1 => n8163, B2 => 
                           n5043, ZN => n8231);
   U9064 : AOI22_X1 port map( A1 => n8164, A2 => n5044, B1 => n8165, B2 => 
                           n5045, ZN => n8230);
   U9065 : NAND3_X1 port map( A1 => n8234, A2 => n8235, A3 => n8236, ZN => 
                           n12494);
   U9066 : AOI221_X1 port map( B1 => n8159, B2 => n5049, C1 => n189, C2 => 
                           MEM_IN(18), A => n8237, ZN => n8236);
   U9067 : OAI22_X1 port map( A1 => n11131, A2 => n287, B1 => n5051, B2 => n138
                           , ZN => n8237);
   U9068 : AOI22_X1 port map( A1 => n8162, A2 => n5052, B1 => n8163, B2 => 
                           n5053, ZN => n8235);
   U9069 : AOI22_X1 port map( A1 => n8164, A2 => n5054, B1 => n8165, B2 => 
                           n5055, ZN => n8234);
   U9070 : NAND3_X1 port map( A1 => n8238, A2 => n8239, A3 => n8240, ZN => 
                           n12493);
   U9071 : AOI221_X1 port map( B1 => n8159, B2 => n5059, C1 => n189, C2 => 
                           MEM_IN(19), A => n8241, ZN => n8240);
   U9072 : OAI22_X1 port map( A1 => n11130, A2 => n287, B1 => n5061, B2 => n138
                           , ZN => n8241);
   U9073 : AOI22_X1 port map( A1 => n8162, A2 => n5062, B1 => n8163, B2 => 
                           n5063, ZN => n8239);
   U9074 : AOI22_X1 port map( A1 => n8164, A2 => n5064, B1 => n8165, B2 => 
                           n5065, ZN => n8238);
   U9075 : NAND3_X1 port map( A1 => n8242, A2 => n8243, A3 => n8244, ZN => 
                           n12492);
   U9076 : AOI221_X1 port map( B1 => n8159, B2 => n5069, C1 => n189, C2 => 
                           MEM_IN(20), A => n8245, ZN => n8244);
   U9077 : OAI22_X1 port map( A1 => n11129, A2 => n287, B1 => n5071, B2 => n138
                           , ZN => n8245);
   U9078 : AOI22_X1 port map( A1 => n8162, A2 => n5072, B1 => n8163, B2 => 
                           n5073, ZN => n8243);
   U9079 : AOI22_X1 port map( A1 => n8164, A2 => n5074, B1 => n8165, B2 => 
                           n5075, ZN => n8242);
   U9080 : NAND3_X1 port map( A1 => n8246, A2 => n8247, A3 => n8248, ZN => 
                           n12491);
   U9081 : AOI221_X1 port map( B1 => n8159, B2 => n5079, C1 => n189, C2 => 
                           MEM_IN(21), A => n8249, ZN => n8248);
   U9082 : OAI22_X1 port map( A1 => n11128, A2 => n287, B1 => n5081, B2 => n138
                           , ZN => n8249);
   U9083 : AOI22_X1 port map( A1 => n8162, A2 => n5082, B1 => n8163, B2 => 
                           n5083, ZN => n8247);
   U9084 : AOI22_X1 port map( A1 => n8164, A2 => n5084, B1 => n8165, B2 => 
                           n5085, ZN => n8246);
   U9085 : NAND3_X1 port map( A1 => n8250, A2 => n8251, A3 => n8252, ZN => 
                           n12490);
   U9086 : AOI221_X1 port map( B1 => n8159, B2 => n5089, C1 => n189, C2 => 
                           MEM_IN(22), A => n8253, ZN => n8252);
   U9087 : OAI22_X1 port map( A1 => n11127, A2 => n287, B1 => n5091, B2 => n138
                           , ZN => n8253);
   U9088 : AOI22_X1 port map( A1 => n8162, A2 => n5092, B1 => n8163, B2 => 
                           n5093, ZN => n8251);
   U9089 : AOI22_X1 port map( A1 => n8164, A2 => n5094, B1 => n8165, B2 => 
                           n5095, ZN => n8250);
   U9090 : NAND3_X1 port map( A1 => n8254, A2 => n8255, A3 => n8256, ZN => 
                           n12489);
   U9091 : AOI221_X1 port map( B1 => n8159, B2 => n5099, C1 => n189, C2 => 
                           MEM_IN(23), A => n8257, ZN => n8256);
   U9092 : OAI22_X1 port map( A1 => n11126, A2 => n287, B1 => n5101, B2 => n138
                           , ZN => n8257);
   U9093 : AOI22_X1 port map( A1 => n8162, A2 => n5102, B1 => n8163, B2 => 
                           n5103, ZN => n8255);
   U9094 : AOI22_X1 port map( A1 => n8164, A2 => n5104, B1 => n8165, B2 => 
                           n5105, ZN => n8254);
   U9095 : NAND3_X1 port map( A1 => n8258, A2 => n8259, A3 => n8260, ZN => 
                           n12488);
   U9096 : AOI221_X1 port map( B1 => n8159, B2 => n5109, C1 => n189, C2 => 
                           MEM_IN(24), A => n8261, ZN => n8260);
   U9097 : OAI22_X1 port map( A1 => n11125, A2 => n287, B1 => n5111, B2 => n138
                           , ZN => n8261);
   U9098 : AOI22_X1 port map( A1 => n8162, A2 => n5112, B1 => n8163, B2 => 
                           n5113, ZN => n8259);
   U9099 : AOI22_X1 port map( A1 => n8164, A2 => n5114, B1 => n8165, B2 => 
                           n5115, ZN => n8258);
   U9100 : NAND3_X1 port map( A1 => n8262, A2 => n8263, A3 => n8264, ZN => 
                           n12487);
   U9101 : AOI221_X1 port map( B1 => n8159, B2 => n5119, C1 => n189, C2 => 
                           MEM_IN(25), A => n8265, ZN => n8264);
   U9102 : OAI22_X1 port map( A1 => n11124, A2 => n287, B1 => n5121, B2 => n138
                           , ZN => n8265);
   U9103 : AOI22_X1 port map( A1 => n8162, A2 => n5122, B1 => n8163, B2 => 
                           n5123, ZN => n8263);
   U9104 : AOI22_X1 port map( A1 => n8164, A2 => n5124, B1 => n8165, B2 => 
                           n5125, ZN => n8262);
   U9105 : NAND3_X1 port map( A1 => n8266, A2 => n8267, A3 => n8268, ZN => 
                           n12486);
   U9106 : AOI221_X1 port map( B1 => n8159, B2 => n5129, C1 => n189, C2 => 
                           MEM_IN(26), A => n8269, ZN => n8268);
   U9107 : OAI22_X1 port map( A1 => n11123, A2 => n287, B1 => n5131, B2 => n138
                           , ZN => n8269);
   U9108 : AOI22_X1 port map( A1 => n8162, A2 => n5132, B1 => n8163, B2 => 
                           n5133, ZN => n8267);
   U9109 : AOI22_X1 port map( A1 => n8164, A2 => n5134, B1 => n8165, B2 => 
                           n5135, ZN => n8266);
   U9110 : NAND3_X1 port map( A1 => n8270, A2 => n8271, A3 => n8272, ZN => 
                           n12485);
   U9111 : AOI221_X1 port map( B1 => n8159, B2 => n5139, C1 => n189, C2 => 
                           MEM_IN(27), A => n8273, ZN => n8272);
   U9112 : OAI22_X1 port map( A1 => n11122, A2 => n287, B1 => n5141, B2 => n138
                           , ZN => n8273);
   U9113 : AOI22_X1 port map( A1 => n8162, A2 => n5142, B1 => n8163, B2 => 
                           n5143, ZN => n8271);
   U9114 : AOI22_X1 port map( A1 => n8164, A2 => n5144, B1 => n8165, B2 => 
                           n5145, ZN => n8270);
   U9115 : NAND3_X1 port map( A1 => n8274, A2 => n8275, A3 => n8276, ZN => 
                           n12484);
   U9116 : AOI221_X1 port map( B1 => n8159, B2 => n5149, C1 => n189, C2 => 
                           MEM_IN(28), A => n8277, ZN => n8276);
   U9117 : OAI22_X1 port map( A1 => n11121, A2 => n287, B1 => n5151, B2 => n138
                           , ZN => n8277);
   U9118 : AOI22_X1 port map( A1 => n8162, A2 => n5152, B1 => n8163, B2 => 
                           n5153, ZN => n8275);
   U9119 : AOI22_X1 port map( A1 => n8164, A2 => n5154, B1 => n8165, B2 => 
                           n5155, ZN => n8274);
   U9120 : NAND3_X1 port map( A1 => n8278, A2 => n8279, A3 => n8280, ZN => 
                           n12483);
   U9121 : AOI221_X1 port map( B1 => n8159, B2 => n5159, C1 => n189, C2 => 
                           MEM_IN(29), A => n8281, ZN => n8280);
   U9122 : OAI22_X1 port map( A1 => n11120, A2 => n287, B1 => n5161, B2 => n138
                           , ZN => n8281);
   U9123 : AOI22_X1 port map( A1 => n8162, A2 => n5162, B1 => n8163, B2 => 
                           n5163, ZN => n8279);
   U9124 : AOI22_X1 port map( A1 => n8164, A2 => n5164, B1 => n8165, B2 => 
                           n5165, ZN => n8278);
   U9125 : NAND3_X1 port map( A1 => n8282, A2 => n8283, A3 => n8284, ZN => 
                           n12482);
   U9126 : AOI221_X1 port map( B1 => n8159, B2 => n5169, C1 => n189, C2 => 
                           MEM_IN(30), A => n8285, ZN => n8284);
   U9127 : OAI22_X1 port map( A1 => n11119, A2 => n287, B1 => n5171, B2 => n138
                           , ZN => n8285);
   U9128 : AOI22_X1 port map( A1 => n8162, A2 => n5172, B1 => n8163, B2 => 
                           n5173, ZN => n8283);
   U9129 : AOI22_X1 port map( A1 => n8164, A2 => n5174, B1 => n8165, B2 => 
                           n5175, ZN => n8282);
   U9130 : NAND3_X1 port map( A1 => n8286, A2 => n8287, A3 => n8288, ZN => 
                           n12481);
   U9131 : AOI221_X1 port map( B1 => n8159, B2 => n5179, C1 => n189, C2 => 
                           MEM_IN(31), A => n8289, ZN => n8288);
   U9132 : OAI22_X1 port map( A1 => n11118, A2 => n287, B1 => n5181, B2 => n138
                           , ZN => n8289);
   U9133 : INV_X1 port map( A => n8293, ZN => n8292);
   U9134 : INV_X1 port map( A => n7850, ZN => n7847);
   U9135 : AOI22_X1 port map( A1 => n8162, A2 => n5191, B1 => n8163, B2 => 
                           n5192, ZN => n8287);
   U9136 : AOI22_X1 port map( A1 => n8164, A2 => n5195, B1 => n8165, B2 => 
                           n5196, ZN => n8286);
   U9137 : OAI22_X1 port map( A1 => n8293, A2 => n8291, B1 => n208, B2 => n286,
                           ZN => n8294);
   U9138 : NAND3_X1 port map( A1 => n208, A2 => n287, A3 => n7265, ZN => n8291)
                           ;
   U9139 : INV_X1 port map( A => n8290, ZN => n7265);
   U9140 : OAI22_X1 port map( A1 => n4786, A2 => n8297, B1 => n8298, B2 => 
                           n5204, ZN => n8161);
   U9141 : NOR2_X1 port map( A1 => n8290, A2 => n8293, ZN => n8298);
   U9142 : NAND3_X1 port map( A1 => n8002, A2 => n7413, A3 => n8299, ZN => 
                           n8290);
   U9143 : AOI211_X1 port map( C1 => n7705, C2 => n8300, A => n8301, B => n7850
                           , ZN => n8297);
   U9144 : NOR2_X1 port map( A1 => n7413, A2 => n4787, ZN => n7850);
   U9145 : INV_X1 port map( A => n5923, ZN => n8300);
   U9146 : NAND2_X1 port map( A1 => n8302, A2 => n8303, ZN => n8293);
   U9147 : NOR2_X1 port map( A1 => n8147, A2 => n7413, ZN => n8146);
   U9148 : NAND2_X1 port map( A1 => n7708, A2 => n5926, ZN => n7413);
   U9149 : NAND3_X1 port map( A1 => n8304, A2 => n8305, A3 => n8306, ZN => 
                           n12480);
   U9150 : AOI221_X1 port map( B1 => n8307, B2 => n4863, C1 => n182, C2 => 
                           MEM_IN(0), A => n8308, ZN => n8306);
   U9151 : OAI22_X1 port map( A1 => n11117, A2 => n289, B1 => n4867, B2 => n139
                           , ZN => n8308);
   U9152 : AOI22_X1 port map( A1 => n8310, A2 => n4869, B1 => n8311, B2 => 
                           n4871, ZN => n8305);
   U9153 : AOI22_X1 port map( A1 => n8312, A2 => n4873, B1 => n8313, B2 => 
                           n4875, ZN => n8304);
   U9154 : NAND3_X1 port map( A1 => n8314, A2 => n8315, A3 => n8316, ZN => 
                           n12479);
   U9155 : AOI221_X1 port map( B1 => n8307, B2 => n4879, C1 => n182, C2 => 
                           MEM_IN(1), A => n8317, ZN => n8316);
   U9156 : OAI22_X1 port map( A1 => n11116, A2 => n289, B1 => n4881, B2 => n139
                           , ZN => n8317);
   U9157 : AOI22_X1 port map( A1 => n8310, A2 => n4882, B1 => n8311, B2 => 
                           n4883, ZN => n8315);
   U9158 : AOI22_X1 port map( A1 => n8312, A2 => n4884, B1 => n8313, B2 => 
                           n4885, ZN => n8314);
   U9159 : NAND3_X1 port map( A1 => n8318, A2 => n8319, A3 => n8320, ZN => 
                           n12478);
   U9160 : AOI221_X1 port map( B1 => n8307, B2 => n4889, C1 => n182, C2 => 
                           MEM_IN(2), A => n8321, ZN => n8320);
   U9161 : OAI22_X1 port map( A1 => n11115, A2 => n289, B1 => n4891, B2 => n139
                           , ZN => n8321);
   U9162 : AOI22_X1 port map( A1 => n8310, A2 => n4892, B1 => n8311, B2 => 
                           n4893, ZN => n8319);
   U9163 : AOI22_X1 port map( A1 => n8312, A2 => n4894, B1 => n8313, B2 => 
                           n4895, ZN => n8318);
   U9164 : NAND3_X1 port map( A1 => n8322, A2 => n8323, A3 => n8324, ZN => 
                           n12477);
   U9165 : AOI221_X1 port map( B1 => n8307, B2 => n4899, C1 => n182, C2 => 
                           MEM_IN(3), A => n8325, ZN => n8324);
   U9166 : OAI22_X1 port map( A1 => n11114, A2 => n289, B1 => n4901, B2 => n139
                           , ZN => n8325);
   U9167 : AOI22_X1 port map( A1 => n8310, A2 => n4902, B1 => n8311, B2 => 
                           n4903, ZN => n8323);
   U9168 : AOI22_X1 port map( A1 => n8312, A2 => n4904, B1 => n8313, B2 => 
                           n4905, ZN => n8322);
   U9169 : NAND3_X1 port map( A1 => n8326, A2 => n8327, A3 => n8328, ZN => 
                           n12476);
   U9170 : AOI221_X1 port map( B1 => n8307, B2 => n4909, C1 => n182, C2 => 
                           MEM_IN(4), A => n8329, ZN => n8328);
   U9171 : OAI22_X1 port map( A1 => n11113, A2 => n289, B1 => n4911, B2 => n139
                           , ZN => n8329);
   U9172 : AOI22_X1 port map( A1 => n8310, A2 => n4912, B1 => n8311, B2 => 
                           n4913, ZN => n8327);
   U9173 : AOI22_X1 port map( A1 => n8312, A2 => n4914, B1 => n8313, B2 => 
                           n4915, ZN => n8326);
   U9174 : NAND3_X1 port map( A1 => n8330, A2 => n8331, A3 => n8332, ZN => 
                           n12475);
   U9175 : AOI221_X1 port map( B1 => n8307, B2 => n4919, C1 => n182, C2 => 
                           MEM_IN(5), A => n8333, ZN => n8332);
   U9176 : OAI22_X1 port map( A1 => n11112, A2 => n289, B1 => n4921, B2 => n139
                           , ZN => n8333);
   U9177 : AOI22_X1 port map( A1 => n8310, A2 => n4922, B1 => n8311, B2 => 
                           n4923, ZN => n8331);
   U9178 : AOI22_X1 port map( A1 => n8312, A2 => n4924, B1 => n8313, B2 => 
                           n4925, ZN => n8330);
   U9179 : NAND3_X1 port map( A1 => n8334, A2 => n8335, A3 => n8336, ZN => 
                           n12474);
   U9180 : AOI221_X1 port map( B1 => n8307, B2 => n4929, C1 => n182, C2 => 
                           MEM_IN(6), A => n8337, ZN => n8336);
   U9181 : OAI22_X1 port map( A1 => n11111, A2 => n289, B1 => n4931, B2 => n139
                           , ZN => n8337);
   U9182 : AOI22_X1 port map( A1 => n8310, A2 => n4932, B1 => n8311, B2 => 
                           n4933, ZN => n8335);
   U9183 : AOI22_X1 port map( A1 => n8312, A2 => n4934, B1 => n8313, B2 => 
                           n4935, ZN => n8334);
   U9184 : NAND3_X1 port map( A1 => n8338, A2 => n8339, A3 => n8340, ZN => 
                           n12473);
   U9185 : AOI221_X1 port map( B1 => n8307, B2 => n4939, C1 => n182, C2 => 
                           MEM_IN(7), A => n8341, ZN => n8340);
   U9186 : OAI22_X1 port map( A1 => n11110, A2 => n289, B1 => n4941, B2 => n139
                           , ZN => n8341);
   U9187 : AOI22_X1 port map( A1 => n8310, A2 => n4942, B1 => n8311, B2 => 
                           n4943, ZN => n8339);
   U9188 : AOI22_X1 port map( A1 => n8312, A2 => n4944, B1 => n8313, B2 => 
                           n4945, ZN => n8338);
   U9189 : NAND3_X1 port map( A1 => n8342, A2 => n8343, A3 => n8344, ZN => 
                           n12472);
   U9190 : AOI221_X1 port map( B1 => n8307, B2 => n4949, C1 => n182, C2 => 
                           MEM_IN(8), A => n8345, ZN => n8344);
   U9191 : OAI22_X1 port map( A1 => n11109, A2 => n289, B1 => n4951, B2 => n139
                           , ZN => n8345);
   U9192 : AOI22_X1 port map( A1 => n8310, A2 => n4952, B1 => n8311, B2 => 
                           n4953, ZN => n8343);
   U9193 : AOI22_X1 port map( A1 => n8312, A2 => n4954, B1 => n8313, B2 => 
                           n4955, ZN => n8342);
   U9194 : NAND3_X1 port map( A1 => n8346, A2 => n8347, A3 => n8348, ZN => 
                           n12471);
   U9195 : AOI221_X1 port map( B1 => n8307, B2 => n4959, C1 => n182, C2 => 
                           MEM_IN(9), A => n8349, ZN => n8348);
   U9196 : OAI22_X1 port map( A1 => n11108, A2 => n289, B1 => n4961, B2 => n139
                           , ZN => n8349);
   U9197 : AOI22_X1 port map( A1 => n8310, A2 => n4962, B1 => n8311, B2 => 
                           n4963, ZN => n8347);
   U9198 : AOI22_X1 port map( A1 => n8312, A2 => n4964, B1 => n8313, B2 => 
                           n4965, ZN => n8346);
   U9199 : NAND3_X1 port map( A1 => n8350, A2 => n8351, A3 => n8352, ZN => 
                           n12470);
   U9200 : AOI221_X1 port map( B1 => n8307, B2 => n4969, C1 => n182, C2 => 
                           MEM_IN(10), A => n8353, ZN => n8352);
   U9201 : OAI22_X1 port map( A1 => n11107, A2 => n289, B1 => n4971, B2 => n139
                           , ZN => n8353);
   U9202 : AOI22_X1 port map( A1 => n8310, A2 => n4972, B1 => n8311, B2 => 
                           n4973, ZN => n8351);
   U9203 : AOI22_X1 port map( A1 => n8312, A2 => n4974, B1 => n8313, B2 => 
                           n4975, ZN => n8350);
   U9204 : NAND3_X1 port map( A1 => n8354, A2 => n8355, A3 => n8356, ZN => 
                           n12469);
   U9205 : AOI221_X1 port map( B1 => n8307, B2 => n4979, C1 => n182, C2 => 
                           MEM_IN(11), A => n8357, ZN => n8356);
   U9206 : OAI22_X1 port map( A1 => n11106, A2 => n289, B1 => n4981, B2 => n139
                           , ZN => n8357);
   U9207 : AOI22_X1 port map( A1 => n8310, A2 => n4982, B1 => n8311, B2 => 
                           n4983, ZN => n8355);
   U9208 : AOI22_X1 port map( A1 => n8312, A2 => n4984, B1 => n8313, B2 => 
                           n4985, ZN => n8354);
   U9209 : NAND3_X1 port map( A1 => n8358, A2 => n8359, A3 => n8360, ZN => 
                           n12468);
   U9210 : AOI221_X1 port map( B1 => n8307, B2 => n4989, C1 => n182, C2 => 
                           MEM_IN(12), A => n8361, ZN => n8360);
   U9211 : OAI22_X1 port map( A1 => n11105, A2 => n289, B1 => n4991, B2 => n139
                           , ZN => n8361);
   U9212 : AOI22_X1 port map( A1 => n8310, A2 => n4992, B1 => n8311, B2 => 
                           n4993, ZN => n8359);
   U9213 : AOI22_X1 port map( A1 => n8312, A2 => n4994, B1 => n8313, B2 => 
                           n4995, ZN => n8358);
   U9214 : NAND3_X1 port map( A1 => n8362, A2 => n8363, A3 => n8364, ZN => 
                           n12467);
   U9215 : AOI221_X1 port map( B1 => n8307, B2 => n4999, C1 => n182, C2 => 
                           MEM_IN(13), A => n8365, ZN => n8364);
   U9216 : OAI22_X1 port map( A1 => n11104, A2 => n289, B1 => n5001, B2 => n139
                           , ZN => n8365);
   U9217 : AOI22_X1 port map( A1 => n8310, A2 => n5002, B1 => n8311, B2 => 
                           n5003, ZN => n8363);
   U9218 : AOI22_X1 port map( A1 => n8312, A2 => n5004, B1 => n8313, B2 => 
                           n5005, ZN => n8362);
   U9219 : NAND3_X1 port map( A1 => n8366, A2 => n8367, A3 => n8368, ZN => 
                           n12466);
   U9220 : AOI221_X1 port map( B1 => n8307, B2 => n5009, C1 => n182, C2 => 
                           MEM_IN(14), A => n8369, ZN => n8368);
   U9221 : OAI22_X1 port map( A1 => n11103, A2 => n289, B1 => n5011, B2 => n139
                           , ZN => n8369);
   U9222 : AOI22_X1 port map( A1 => n8310, A2 => n5012, B1 => n8311, B2 => 
                           n5013, ZN => n8367);
   U9223 : AOI22_X1 port map( A1 => n8312, A2 => n5014, B1 => n8313, B2 => 
                           n5015, ZN => n8366);
   U9224 : NAND3_X1 port map( A1 => n8370, A2 => n8371, A3 => n8372, ZN => 
                           n12465);
   U9225 : AOI221_X1 port map( B1 => n8307, B2 => n5019, C1 => n182, C2 => 
                           MEM_IN(15), A => n8373, ZN => n8372);
   U9226 : OAI22_X1 port map( A1 => n11102, A2 => n289, B1 => n5021, B2 => n139
                           , ZN => n8373);
   U9227 : AOI22_X1 port map( A1 => n8310, A2 => n5022, B1 => n8311, B2 => 
                           n5023, ZN => n8371);
   U9228 : AOI22_X1 port map( A1 => n8312, A2 => n5024, B1 => n8313, B2 => 
                           n5025, ZN => n8370);
   U9229 : NAND3_X1 port map( A1 => n8374, A2 => n8375, A3 => n8376, ZN => 
                           n12464);
   U9230 : AOI221_X1 port map( B1 => n8307, B2 => n5029, C1 => n182, C2 => 
                           MEM_IN(16), A => n8377, ZN => n8376);
   U9231 : OAI22_X1 port map( A1 => n11101, A2 => n289, B1 => n5031, B2 => n139
                           , ZN => n8377);
   U9232 : AOI22_X1 port map( A1 => n8310, A2 => n5032, B1 => n8311, B2 => 
                           n5033, ZN => n8375);
   U9233 : AOI22_X1 port map( A1 => n8312, A2 => n5034, B1 => n8313, B2 => 
                           n5035, ZN => n8374);
   U9234 : NAND3_X1 port map( A1 => n8378, A2 => n8379, A3 => n8380, ZN => 
                           n12463);
   U9235 : AOI221_X1 port map( B1 => n8307, B2 => n5039, C1 => n182, C2 => 
                           MEM_IN(17), A => n8381, ZN => n8380);
   U9236 : OAI22_X1 port map( A1 => n11100, A2 => n289, B1 => n5041, B2 => n139
                           , ZN => n8381);
   U9237 : AOI22_X1 port map( A1 => n8310, A2 => n5042, B1 => n8311, B2 => 
                           n5043, ZN => n8379);
   U9238 : AOI22_X1 port map( A1 => n8312, A2 => n5044, B1 => n8313, B2 => 
                           n5045, ZN => n8378);
   U9239 : NAND3_X1 port map( A1 => n8382, A2 => n8383, A3 => n8384, ZN => 
                           n12462);
   U9240 : AOI221_X1 port map( B1 => n8307, B2 => n5049, C1 => n182, C2 => 
                           MEM_IN(18), A => n8385, ZN => n8384);
   U9241 : OAI22_X1 port map( A1 => n11099, A2 => n289, B1 => n5051, B2 => n139
                           , ZN => n8385);
   U9242 : AOI22_X1 port map( A1 => n8310, A2 => n5052, B1 => n8311, B2 => 
                           n5053, ZN => n8383);
   U9243 : AOI22_X1 port map( A1 => n8312, A2 => n5054, B1 => n8313, B2 => 
                           n5055, ZN => n8382);
   U9244 : NAND3_X1 port map( A1 => n8386, A2 => n8387, A3 => n8388, ZN => 
                           n12461);
   U9245 : AOI221_X1 port map( B1 => n8307, B2 => n5059, C1 => n182, C2 => 
                           MEM_IN(19), A => n8389, ZN => n8388);
   U9246 : OAI22_X1 port map( A1 => n11098, A2 => n289, B1 => n5061, B2 => n139
                           , ZN => n8389);
   U9247 : AOI22_X1 port map( A1 => n8310, A2 => n5062, B1 => n8311, B2 => 
                           n5063, ZN => n8387);
   U9248 : AOI22_X1 port map( A1 => n8312, A2 => n5064, B1 => n8313, B2 => 
                           n5065, ZN => n8386);
   U9249 : NAND3_X1 port map( A1 => n8390, A2 => n8391, A3 => n8392, ZN => 
                           n12460);
   U9250 : AOI221_X1 port map( B1 => n8307, B2 => n5069, C1 => n182, C2 => 
                           MEM_IN(20), A => n8393, ZN => n8392);
   U9251 : OAI22_X1 port map( A1 => n11097, A2 => n289, B1 => n5071, B2 => n139
                           , ZN => n8393);
   U9252 : AOI22_X1 port map( A1 => n8310, A2 => n5072, B1 => n8311, B2 => 
                           n5073, ZN => n8391);
   U9253 : AOI22_X1 port map( A1 => n8312, A2 => n5074, B1 => n8313, B2 => 
                           n5075, ZN => n8390);
   U9254 : NAND3_X1 port map( A1 => n8394, A2 => n8395, A3 => n8396, ZN => 
                           n12459);
   U9255 : AOI221_X1 port map( B1 => n8307, B2 => n5079, C1 => n182, C2 => 
                           MEM_IN(21), A => n8397, ZN => n8396);
   U9256 : OAI22_X1 port map( A1 => n11096, A2 => n289, B1 => n5081, B2 => n139
                           , ZN => n8397);
   U9257 : AOI22_X1 port map( A1 => n8310, A2 => n5082, B1 => n8311, B2 => 
                           n5083, ZN => n8395);
   U9258 : AOI22_X1 port map( A1 => n8312, A2 => n5084, B1 => n8313, B2 => 
                           n5085, ZN => n8394);
   U9259 : NAND3_X1 port map( A1 => n8398, A2 => n8399, A3 => n8400, ZN => 
                           n12458);
   U9260 : AOI221_X1 port map( B1 => n8307, B2 => n5089, C1 => n182, C2 => 
                           MEM_IN(22), A => n8401, ZN => n8400);
   U9261 : OAI22_X1 port map( A1 => n11095, A2 => n289, B1 => n5091, B2 => n139
                           , ZN => n8401);
   U9262 : AOI22_X1 port map( A1 => n8310, A2 => n5092, B1 => n8311, B2 => 
                           n5093, ZN => n8399);
   U9263 : AOI22_X1 port map( A1 => n8312, A2 => n5094, B1 => n8313, B2 => 
                           n5095, ZN => n8398);
   U9264 : NAND3_X1 port map( A1 => n8402, A2 => n8403, A3 => n8404, ZN => 
                           n12457);
   U9265 : AOI221_X1 port map( B1 => n8307, B2 => n5099, C1 => n182, C2 => 
                           MEM_IN(23), A => n8405, ZN => n8404);
   U9266 : OAI22_X1 port map( A1 => n11094, A2 => n289, B1 => n5101, B2 => n139
                           , ZN => n8405);
   U9267 : AOI22_X1 port map( A1 => n8310, A2 => n5102, B1 => n8311, B2 => 
                           n5103, ZN => n8403);
   U9268 : AOI22_X1 port map( A1 => n8312, A2 => n5104, B1 => n8313, B2 => 
                           n5105, ZN => n8402);
   U9269 : NAND3_X1 port map( A1 => n8406, A2 => n8407, A3 => n8408, ZN => 
                           n12456);
   U9270 : AOI221_X1 port map( B1 => n8307, B2 => n5109, C1 => n182, C2 => 
                           MEM_IN(24), A => n8409, ZN => n8408);
   U9271 : OAI22_X1 port map( A1 => n11093, A2 => n289, B1 => n5111, B2 => n139
                           , ZN => n8409);
   U9272 : AOI22_X1 port map( A1 => n8310, A2 => n5112, B1 => n8311, B2 => 
                           n5113, ZN => n8407);
   U9273 : AOI22_X1 port map( A1 => n8312, A2 => n5114, B1 => n8313, B2 => 
                           n5115, ZN => n8406);
   U9274 : NAND3_X1 port map( A1 => n8410, A2 => n8411, A3 => n8412, ZN => 
                           n12455);
   U9275 : AOI221_X1 port map( B1 => n8307, B2 => n5119, C1 => n182, C2 => 
                           MEM_IN(25), A => n8413, ZN => n8412);
   U9276 : OAI22_X1 port map( A1 => n11092, A2 => n289, B1 => n5121, B2 => n139
                           , ZN => n8413);
   U9277 : AOI22_X1 port map( A1 => n8310, A2 => n5122, B1 => n8311, B2 => 
                           n5123, ZN => n8411);
   U9278 : AOI22_X1 port map( A1 => n8312, A2 => n5124, B1 => n8313, B2 => 
                           n5125, ZN => n8410);
   U9279 : NAND3_X1 port map( A1 => n8414, A2 => n8415, A3 => n8416, ZN => 
                           n12454);
   U9280 : AOI221_X1 port map( B1 => n8307, B2 => n5129, C1 => n182, C2 => 
                           MEM_IN(26), A => n8417, ZN => n8416);
   U9281 : OAI22_X1 port map( A1 => n11091, A2 => n289, B1 => n5131, B2 => n139
                           , ZN => n8417);
   U9282 : AOI22_X1 port map( A1 => n8310, A2 => n5132, B1 => n8311, B2 => 
                           n5133, ZN => n8415);
   U9283 : AOI22_X1 port map( A1 => n8312, A2 => n5134, B1 => n8313, B2 => 
                           n5135, ZN => n8414);
   U9284 : NAND3_X1 port map( A1 => n8418, A2 => n8419, A3 => n8420, ZN => 
                           n12453);
   U9285 : AOI221_X1 port map( B1 => n8307, B2 => n5139, C1 => n182, C2 => 
                           MEM_IN(27), A => n8421, ZN => n8420);
   U9286 : OAI22_X1 port map( A1 => n11090, A2 => n289, B1 => n5141, B2 => n139
                           , ZN => n8421);
   U9287 : AOI22_X1 port map( A1 => n8310, A2 => n5142, B1 => n8311, B2 => 
                           n5143, ZN => n8419);
   U9288 : AOI22_X1 port map( A1 => n8312, A2 => n5144, B1 => n8313, B2 => 
                           n5145, ZN => n8418);
   U9289 : NAND3_X1 port map( A1 => n8422, A2 => n8423, A3 => n8424, ZN => 
                           n12452);
   U9290 : AOI221_X1 port map( B1 => n8307, B2 => n5149, C1 => n182, C2 => 
                           MEM_IN(28), A => n8425, ZN => n8424);
   U9291 : OAI22_X1 port map( A1 => n11089, A2 => n289, B1 => n5151, B2 => n139
                           , ZN => n8425);
   U9292 : AOI22_X1 port map( A1 => n8310, A2 => n5152, B1 => n8311, B2 => 
                           n5153, ZN => n8423);
   U9293 : AOI22_X1 port map( A1 => n8312, A2 => n5154, B1 => n8313, B2 => 
                           n5155, ZN => n8422);
   U9294 : NAND3_X1 port map( A1 => n8426, A2 => n8427, A3 => n8428, ZN => 
                           n12451);
   U9295 : AOI221_X1 port map( B1 => n8307, B2 => n5159, C1 => n182, C2 => 
                           MEM_IN(29), A => n8429, ZN => n8428);
   U9296 : OAI22_X1 port map( A1 => n11088, A2 => n289, B1 => n5161, B2 => n139
                           , ZN => n8429);
   U9297 : AOI22_X1 port map( A1 => n8310, A2 => n5162, B1 => n8311, B2 => 
                           n5163, ZN => n8427);
   U9298 : AOI22_X1 port map( A1 => n8312, A2 => n5164, B1 => n8313, B2 => 
                           n5165, ZN => n8426);
   U9299 : NAND3_X1 port map( A1 => n8430, A2 => n8431, A3 => n8432, ZN => 
                           n12450);
   U9300 : AOI221_X1 port map( B1 => n8307, B2 => n5169, C1 => n182, C2 => 
                           MEM_IN(30), A => n8433, ZN => n8432);
   U9301 : OAI22_X1 port map( A1 => n11087, A2 => n289, B1 => n5171, B2 => n139
                           , ZN => n8433);
   U9302 : AOI22_X1 port map( A1 => n8310, A2 => n5172, B1 => n8311, B2 => 
                           n5173, ZN => n8431);
   U9303 : AOI22_X1 port map( A1 => n8312, A2 => n5174, B1 => n8313, B2 => 
                           n5175, ZN => n8430);
   U9304 : NAND3_X1 port map( A1 => n8434, A2 => n8435, A3 => n8436, ZN => 
                           n12449);
   U9305 : AOI221_X1 port map( B1 => n8307, B2 => n5179, C1 => n182, C2 => 
                           MEM_IN(31), A => n8437, ZN => n8436);
   U9306 : OAI22_X1 port map( A1 => n11086, A2 => n289, B1 => n5181, B2 => n139
                           , ZN => n8437);
   U9307 : INV_X1 port map( A => n8441, ZN => n8440);
   U9308 : NAND2_X1 port map( A1 => n5206, A2 => n8147, ZN => n8142);
   U9309 : NAND2_X1 port map( A1 => n7853, A2 => n5206, ZN => n8147);
   U9310 : AOI22_X1 port map( A1 => n8310, A2 => n5191, B1 => n8311, B2 => 
                           n5192, ZN => n8435);
   U9311 : AOI22_X1 port map( A1 => n8312, A2 => n5195, B1 => n8313, B2 => 
                           n5196, ZN => n8434);
   U9312 : OAI22_X1 port map( A1 => n8441, A2 => n8439, B1 => n208, B2 => n288,
                           ZN => n8442);
   U9313 : NAND3_X1 port map( A1 => n208, A2 => n289, A3 => n7412, ZN => n8439)
                           ;
   U9314 : INV_X1 port map( A => n8438, ZN => n7412);
   U9315 : OAI22_X1 port map( A1 => n4786, A2 => n8445, B1 => n8446, B2 => 
                           n5204, ZN => n8309);
   U9316 : NOR2_X1 port map( A1 => n8438, A2 => n8441, ZN => n8446);
   U9317 : NAND2_X1 port map( A1 => n8447, A2 => n8002, ZN => n8438);
   U9318 : AOI211_X1 port map( C1 => n7705, C2 => n8448, A => n8301, B => n8444
                           , ZN => n8445);
   U9319 : OAI21_X1 port map( B1 => n8002, B2 => n4787, A => n5368, ZN => n8301
                           );
   U9320 : AND2_X1 port map( A1 => n7853, A2 => n7858, ZN => n8002);
   U9321 : AND2_X1 port map( A1 => n7707, A2 => n7562, ZN => n7853);
   U9322 : INV_X1 port map( A => n7856, ZN => n7705);
   U9323 : NAND2_X1 port map( A1 => n8449, A2 => n8450, ZN => n8441);
   U9324 : NOR2_X1 port map( A1 => n7562, A2 => n4787, ZN => n7998);
   U9325 : NAND2_X1 port map( A1 => n7708, A2 => n6079, ZN => n7562);
   U9326 : NAND3_X1 port map( A1 => n8451, A2 => n8452, A3 => n8453, ZN => 
                           n12448);
   U9327 : AOI221_X1 port map( B1 => n211, B2 => n4863, C1 => n183, C2 => 
                           MEM_IN(0), A => n8454, ZN => n8453);
   U9328 : OAI22_X1 port map( A1 => n11085, A2 => n267, B1 => n4867, B2 => n136
                           , ZN => n8454);
   U9329 : AOI22_X1 port map( A1 => n201, A2 => n4869, B1 => n159, B2 => n4871,
                           ZN => n8452);
   U9330 : AOI22_X1 port map( A1 => n243, A2 => n4873, B1 => n156, B2 => n4875,
                           ZN => n8451);
   U9331 : NAND3_X1 port map( A1 => n8456, A2 => n8457, A3 => n8458, ZN => 
                           n12447);
   U9332 : AOI221_X1 port map( B1 => n211, B2 => n4879, C1 => n183, C2 => 
                           MEM_IN(1), A => n8459, ZN => n8458);
   U9333 : OAI22_X1 port map( A1 => n11084, A2 => n267, B1 => n4881, B2 => n136
                           , ZN => n8459);
   U9334 : AOI22_X1 port map( A1 => n201, A2 => n4882, B1 => n159, B2 => n4883,
                           ZN => n8457);
   U9335 : AOI22_X1 port map( A1 => n243, A2 => n4884, B1 => n156, B2 => n4885,
                           ZN => n8456);
   U9336 : NAND3_X1 port map( A1 => n8460, A2 => n8461, A3 => n8462, ZN => 
                           n12446);
   U9337 : AOI221_X1 port map( B1 => n211, B2 => n4889, C1 => n183, C2 => 
                           MEM_IN(2), A => n8463, ZN => n8462);
   U9338 : OAI22_X1 port map( A1 => n11083, A2 => n267, B1 => n4891, B2 => n136
                           , ZN => n8463);
   U9339 : AOI22_X1 port map( A1 => n201, A2 => n4892, B1 => n159, B2 => n4893,
                           ZN => n8461);
   U9340 : AOI22_X1 port map( A1 => n243, A2 => n4894, B1 => n156, B2 => n4895,
                           ZN => n8460);
   U9341 : NAND3_X1 port map( A1 => n8464, A2 => n8465, A3 => n8466, ZN => 
                           n12445);
   U9342 : AOI221_X1 port map( B1 => n211, B2 => n4899, C1 => n183, C2 => 
                           MEM_IN(3), A => n8467, ZN => n8466);
   U9343 : OAI22_X1 port map( A1 => n11082, A2 => n267, B1 => n4901, B2 => n136
                           , ZN => n8467);
   U9344 : AOI22_X1 port map( A1 => n201, A2 => n4902, B1 => n159, B2 => n4903,
                           ZN => n8465);
   U9345 : AOI22_X1 port map( A1 => n243, A2 => n4904, B1 => n156, B2 => n4905,
                           ZN => n8464);
   U9346 : NAND3_X1 port map( A1 => n8468, A2 => n8469, A3 => n8470, ZN => 
                           n12444);
   U9347 : AOI221_X1 port map( B1 => n211, B2 => n4909, C1 => n183, C2 => 
                           MEM_IN(4), A => n8471, ZN => n8470);
   U9348 : OAI22_X1 port map( A1 => n11081, A2 => n267, B1 => n4911, B2 => n136
                           , ZN => n8471);
   U9349 : AOI22_X1 port map( A1 => n201, A2 => n4912, B1 => n159, B2 => n4913,
                           ZN => n8469);
   U9350 : AOI22_X1 port map( A1 => n243, A2 => n4914, B1 => n156, B2 => n4915,
                           ZN => n8468);
   U9351 : NAND3_X1 port map( A1 => n8472, A2 => n8473, A3 => n8474, ZN => 
                           n12443);
   U9352 : AOI221_X1 port map( B1 => n211, B2 => n4919, C1 => n183, C2 => 
                           MEM_IN(5), A => n8475, ZN => n8474);
   U9353 : OAI22_X1 port map( A1 => n11080, A2 => n267, B1 => n4921, B2 => n136
                           , ZN => n8475);
   U9354 : AOI22_X1 port map( A1 => n201, A2 => n4922, B1 => n159, B2 => n4923,
                           ZN => n8473);
   U9355 : AOI22_X1 port map( A1 => n243, A2 => n4924, B1 => n156, B2 => n4925,
                           ZN => n8472);
   U9356 : NAND3_X1 port map( A1 => n8476, A2 => n8477, A3 => n8478, ZN => 
                           n12442);
   U9357 : AOI221_X1 port map( B1 => n211, B2 => n4929, C1 => n183, C2 => 
                           MEM_IN(6), A => n8479, ZN => n8478);
   U9358 : OAI22_X1 port map( A1 => n11079, A2 => n267, B1 => n4931, B2 => n136
                           , ZN => n8479);
   U9359 : AOI22_X1 port map( A1 => n201, A2 => n4932, B1 => n159, B2 => n4933,
                           ZN => n8477);
   U9360 : AOI22_X1 port map( A1 => n243, A2 => n4934, B1 => n156, B2 => n4935,
                           ZN => n8476);
   U9361 : NAND3_X1 port map( A1 => n8480, A2 => n8481, A3 => n8482, ZN => 
                           n12441);
   U9362 : AOI221_X1 port map( B1 => n211, B2 => n4939, C1 => n183, C2 => 
                           MEM_IN(7), A => n8483, ZN => n8482);
   U9363 : OAI22_X1 port map( A1 => n11078, A2 => n267, B1 => n4941, B2 => n136
                           , ZN => n8483);
   U9364 : AOI22_X1 port map( A1 => n201, A2 => n4942, B1 => n159, B2 => n4943,
                           ZN => n8481);
   U9365 : AOI22_X1 port map( A1 => n243, A2 => n4944, B1 => n156, B2 => n4945,
                           ZN => n8480);
   U9366 : NAND3_X1 port map( A1 => n8484, A2 => n8485, A3 => n8486, ZN => 
                           n12440);
   U9367 : AOI221_X1 port map( B1 => n211, B2 => n4949, C1 => n183, C2 => 
                           MEM_IN(8), A => n8487, ZN => n8486);
   U9368 : OAI22_X1 port map( A1 => n11077, A2 => n267, B1 => n4951, B2 => n136
                           , ZN => n8487);
   U9369 : AOI22_X1 port map( A1 => n201, A2 => n4952, B1 => n159, B2 => n4953,
                           ZN => n8485);
   U9370 : AOI22_X1 port map( A1 => n243, A2 => n4954, B1 => n156, B2 => n4955,
                           ZN => n8484);
   U9371 : NAND3_X1 port map( A1 => n8488, A2 => n8489, A3 => n8490, ZN => 
                           n12439);
   U9372 : AOI221_X1 port map( B1 => n211, B2 => n4959, C1 => n183, C2 => 
                           MEM_IN(9), A => n8491, ZN => n8490);
   U9373 : OAI22_X1 port map( A1 => n11076, A2 => n267, B1 => n4961, B2 => n136
                           , ZN => n8491);
   U9374 : AOI22_X1 port map( A1 => n201, A2 => n4962, B1 => n159, B2 => n4963,
                           ZN => n8489);
   U9375 : AOI22_X1 port map( A1 => n243, A2 => n4964, B1 => n156, B2 => n4965,
                           ZN => n8488);
   U9376 : NAND3_X1 port map( A1 => n8492, A2 => n8493, A3 => n8494, ZN => 
                           n12438);
   U9377 : AOI221_X1 port map( B1 => n211, B2 => n4969, C1 => n183, C2 => 
                           MEM_IN(10), A => n8495, ZN => n8494);
   U9378 : OAI22_X1 port map( A1 => n11075, A2 => n267, B1 => n4971, B2 => n136
                           , ZN => n8495);
   U9379 : AOI22_X1 port map( A1 => n201, A2 => n4972, B1 => n159, B2 => n4973,
                           ZN => n8493);
   U9380 : AOI22_X1 port map( A1 => n243, A2 => n4974, B1 => n156, B2 => n4975,
                           ZN => n8492);
   U9381 : NAND3_X1 port map( A1 => n8496, A2 => n8497, A3 => n8498, ZN => 
                           n12437);
   U9382 : AOI221_X1 port map( B1 => n211, B2 => n4979, C1 => n183, C2 => 
                           MEM_IN(11), A => n8499, ZN => n8498);
   U9383 : OAI22_X1 port map( A1 => n11074, A2 => n267, B1 => n4981, B2 => n136
                           , ZN => n8499);
   U9384 : AOI22_X1 port map( A1 => n201, A2 => n4982, B1 => n159, B2 => n4983,
                           ZN => n8497);
   U9385 : AOI22_X1 port map( A1 => n243, A2 => n4984, B1 => n156, B2 => n4985,
                           ZN => n8496);
   U9386 : NAND3_X1 port map( A1 => n8500, A2 => n8501, A3 => n8502, ZN => 
                           n12436);
   U9387 : AOI221_X1 port map( B1 => n211, B2 => n4989, C1 => n183, C2 => 
                           MEM_IN(12), A => n8503, ZN => n8502);
   U9388 : OAI22_X1 port map( A1 => n11073, A2 => n267, B1 => n4991, B2 => n136
                           , ZN => n8503);
   U9389 : AOI22_X1 port map( A1 => n201, A2 => n4992, B1 => n159, B2 => n4993,
                           ZN => n8501);
   U9390 : AOI22_X1 port map( A1 => n243, A2 => n4994, B1 => n156, B2 => n4995,
                           ZN => n8500);
   U9391 : NAND3_X1 port map( A1 => n8504, A2 => n8505, A3 => n8506, ZN => 
                           n12435);
   U9392 : AOI221_X1 port map( B1 => n211, B2 => n4999, C1 => n183, C2 => 
                           MEM_IN(13), A => n8507, ZN => n8506);
   U9393 : OAI22_X1 port map( A1 => n11072, A2 => n267, B1 => n5001, B2 => n136
                           , ZN => n8507);
   U9394 : AOI22_X1 port map( A1 => n201, A2 => n5002, B1 => n159, B2 => n5003,
                           ZN => n8505);
   U9395 : AOI22_X1 port map( A1 => n243, A2 => n5004, B1 => n156, B2 => n5005,
                           ZN => n8504);
   U9396 : NAND3_X1 port map( A1 => n8508, A2 => n8509, A3 => n8510, ZN => 
                           n12434);
   U9397 : AOI221_X1 port map( B1 => n211, B2 => n5009, C1 => n183, C2 => 
                           MEM_IN(14), A => n8511, ZN => n8510);
   U9398 : OAI22_X1 port map( A1 => n11071, A2 => n267, B1 => n5011, B2 => n136
                           , ZN => n8511);
   U9399 : AOI22_X1 port map( A1 => n201, A2 => n5012, B1 => n159, B2 => n5013,
                           ZN => n8509);
   U9400 : AOI22_X1 port map( A1 => n243, A2 => n5014, B1 => n156, B2 => n5015,
                           ZN => n8508);
   U9401 : NAND3_X1 port map( A1 => n8512, A2 => n8513, A3 => n8514, ZN => 
                           n12433);
   U9402 : AOI221_X1 port map( B1 => n211, B2 => n5019, C1 => n183, C2 => 
                           MEM_IN(15), A => n8515, ZN => n8514);
   U9403 : OAI22_X1 port map( A1 => n11070, A2 => n267, B1 => n5021, B2 => n136
                           , ZN => n8515);
   U9404 : AOI22_X1 port map( A1 => n201, A2 => n5022, B1 => n159, B2 => n5023,
                           ZN => n8513);
   U9405 : AOI22_X1 port map( A1 => n243, A2 => n5024, B1 => n156, B2 => n5025,
                           ZN => n8512);
   U9406 : NAND3_X1 port map( A1 => n8516, A2 => n8517, A3 => n8518, ZN => 
                           n12432);
   U9407 : AOI221_X1 port map( B1 => n211, B2 => n5029, C1 => n183, C2 => 
                           MEM_IN(16), A => n8519, ZN => n8518);
   U9408 : OAI22_X1 port map( A1 => n11069, A2 => n267, B1 => n5031, B2 => n136
                           , ZN => n8519);
   U9409 : AOI22_X1 port map( A1 => n201, A2 => n5032, B1 => n159, B2 => n5033,
                           ZN => n8517);
   U9410 : AOI22_X1 port map( A1 => n243, A2 => n5034, B1 => n156, B2 => n5035,
                           ZN => n8516);
   U9411 : NAND3_X1 port map( A1 => n8520, A2 => n8521, A3 => n8522, ZN => 
                           n12431);
   U9412 : AOI221_X1 port map( B1 => n211, B2 => n5039, C1 => n183, C2 => 
                           MEM_IN(17), A => n8523, ZN => n8522);
   U9413 : OAI22_X1 port map( A1 => n11068, A2 => n267, B1 => n5041, B2 => n136
                           , ZN => n8523);
   U9414 : AOI22_X1 port map( A1 => n201, A2 => n5042, B1 => n159, B2 => n5043,
                           ZN => n8521);
   U9415 : AOI22_X1 port map( A1 => n243, A2 => n5044, B1 => n156, B2 => n5045,
                           ZN => n8520);
   U9416 : NAND3_X1 port map( A1 => n8524, A2 => n8525, A3 => n8526, ZN => 
                           n12430);
   U9417 : AOI221_X1 port map( B1 => n211, B2 => n5049, C1 => n183, C2 => 
                           MEM_IN(18), A => n8527, ZN => n8526);
   U9418 : OAI22_X1 port map( A1 => n11067, A2 => n267, B1 => n5051, B2 => n136
                           , ZN => n8527);
   U9419 : AOI22_X1 port map( A1 => n201, A2 => n5052, B1 => n159, B2 => n5053,
                           ZN => n8525);
   U9420 : AOI22_X1 port map( A1 => n243, A2 => n5054, B1 => n156, B2 => n5055,
                           ZN => n8524);
   U9421 : NAND3_X1 port map( A1 => n8528, A2 => n8529, A3 => n8530, ZN => 
                           n12429);
   U9422 : AOI221_X1 port map( B1 => n211, B2 => n5059, C1 => n183, C2 => 
                           MEM_IN(19), A => n8531, ZN => n8530);
   U9423 : OAI22_X1 port map( A1 => n11066, A2 => n267, B1 => n5061, B2 => n136
                           , ZN => n8531);
   U9424 : AOI22_X1 port map( A1 => n201, A2 => n5062, B1 => n159, B2 => n5063,
                           ZN => n8529);
   U9425 : AOI22_X1 port map( A1 => n243, A2 => n5064, B1 => n156, B2 => n5065,
                           ZN => n8528);
   U9426 : NAND3_X1 port map( A1 => n8532, A2 => n8533, A3 => n8534, ZN => 
                           n12428);
   U9427 : AOI221_X1 port map( B1 => n211, B2 => n5069, C1 => n183, C2 => 
                           MEM_IN(20), A => n8535, ZN => n8534);
   U9428 : OAI22_X1 port map( A1 => n11065, A2 => n267, B1 => n5071, B2 => n136
                           , ZN => n8535);
   U9429 : AOI22_X1 port map( A1 => n201, A2 => n5072, B1 => n159, B2 => n5073,
                           ZN => n8533);
   U9430 : AOI22_X1 port map( A1 => n243, A2 => n5074, B1 => n156, B2 => n5075,
                           ZN => n8532);
   U9431 : NAND3_X1 port map( A1 => n8536, A2 => n8537, A3 => n8538, ZN => 
                           n12427);
   U9432 : AOI221_X1 port map( B1 => n211, B2 => n5079, C1 => n183, C2 => 
                           MEM_IN(21), A => n8539, ZN => n8538);
   U9433 : OAI22_X1 port map( A1 => n11064, A2 => n267, B1 => n5081, B2 => n136
                           , ZN => n8539);
   U9434 : AOI22_X1 port map( A1 => n201, A2 => n5082, B1 => n159, B2 => n5083,
                           ZN => n8537);
   U9435 : AOI22_X1 port map( A1 => n243, A2 => n5084, B1 => n156, B2 => n5085,
                           ZN => n8536);
   U9436 : NAND3_X1 port map( A1 => n8540, A2 => n8541, A3 => n8542, ZN => 
                           n12426);
   U9437 : AOI221_X1 port map( B1 => n211, B2 => n5089, C1 => n183, C2 => 
                           MEM_IN(22), A => n8543, ZN => n8542);
   U9438 : OAI22_X1 port map( A1 => n11063, A2 => n267, B1 => n5091, B2 => n136
                           , ZN => n8543);
   U9439 : AOI22_X1 port map( A1 => n201, A2 => n5092, B1 => n159, B2 => n5093,
                           ZN => n8541);
   U9440 : AOI22_X1 port map( A1 => n243, A2 => n5094, B1 => n156, B2 => n5095,
                           ZN => n8540);
   U9441 : NAND3_X1 port map( A1 => n8544, A2 => n8545, A3 => n8546, ZN => 
                           n12425);
   U9442 : AOI221_X1 port map( B1 => n211, B2 => n5099, C1 => n183, C2 => 
                           MEM_IN(23), A => n8547, ZN => n8546);
   U9443 : OAI22_X1 port map( A1 => n11062, A2 => n267, B1 => n5101, B2 => n136
                           , ZN => n8547);
   U9444 : AOI22_X1 port map( A1 => n201, A2 => n5102, B1 => n159, B2 => n5103,
                           ZN => n8545);
   U9445 : AOI22_X1 port map( A1 => n243, A2 => n5104, B1 => n156, B2 => n5105,
                           ZN => n8544);
   U9446 : NAND3_X1 port map( A1 => n8548, A2 => n8549, A3 => n8550, ZN => 
                           n12424);
   U9447 : AOI221_X1 port map( B1 => n211, B2 => n5109, C1 => n183, C2 => 
                           MEM_IN(24), A => n8551, ZN => n8550);
   U9448 : OAI22_X1 port map( A1 => n11061, A2 => n267, B1 => n5111, B2 => n136
                           , ZN => n8551);
   U9449 : AOI22_X1 port map( A1 => n201, A2 => n5112, B1 => n159, B2 => n5113,
                           ZN => n8549);
   U9450 : AOI22_X1 port map( A1 => n243, A2 => n5114, B1 => n156, B2 => n5115,
                           ZN => n8548);
   U9451 : NAND3_X1 port map( A1 => n8552, A2 => n8553, A3 => n8554, ZN => 
                           n12423);
   U9452 : AOI221_X1 port map( B1 => n211, B2 => n5119, C1 => n183, C2 => 
                           MEM_IN(25), A => n8555, ZN => n8554);
   U9453 : OAI22_X1 port map( A1 => n11060, A2 => n267, B1 => n5121, B2 => n136
                           , ZN => n8555);
   U9454 : AOI22_X1 port map( A1 => n201, A2 => n5122, B1 => n159, B2 => n5123,
                           ZN => n8553);
   U9455 : AOI22_X1 port map( A1 => n243, A2 => n5124, B1 => n156, B2 => n5125,
                           ZN => n8552);
   U9456 : NAND3_X1 port map( A1 => n8556, A2 => n8557, A3 => n8558, ZN => 
                           n12422);
   U9457 : AOI221_X1 port map( B1 => n211, B2 => n5129, C1 => n183, C2 => 
                           MEM_IN(26), A => n8559, ZN => n8558);
   U9458 : OAI22_X1 port map( A1 => n11059, A2 => n267, B1 => n5131, B2 => n136
                           , ZN => n8559);
   U9459 : AOI22_X1 port map( A1 => n201, A2 => n5132, B1 => n159, B2 => n5133,
                           ZN => n8557);
   U9460 : AOI22_X1 port map( A1 => n243, A2 => n5134, B1 => n156, B2 => n5135,
                           ZN => n8556);
   U9461 : NAND3_X1 port map( A1 => n8560, A2 => n8561, A3 => n8562, ZN => 
                           n12421);
   U9462 : AOI221_X1 port map( B1 => n211, B2 => n5139, C1 => n183, C2 => 
                           MEM_IN(27), A => n8563, ZN => n8562);
   U9463 : OAI22_X1 port map( A1 => n11058, A2 => n267, B1 => n5141, B2 => n136
                           , ZN => n8563);
   U9464 : AOI22_X1 port map( A1 => n201, A2 => n5142, B1 => n159, B2 => n5143,
                           ZN => n8561);
   U9465 : AOI22_X1 port map( A1 => n243, A2 => n5144, B1 => n156, B2 => n5145,
                           ZN => n8560);
   U9466 : NAND3_X1 port map( A1 => n8564, A2 => n8565, A3 => n8566, ZN => 
                           n12420);
   U9467 : AOI221_X1 port map( B1 => n211, B2 => n5149, C1 => n183, C2 => 
                           MEM_IN(28), A => n8567, ZN => n8566);
   U9468 : OAI22_X1 port map( A1 => n11057, A2 => n267, B1 => n5151, B2 => n136
                           , ZN => n8567);
   U9469 : AOI22_X1 port map( A1 => n201, A2 => n5152, B1 => n159, B2 => n5153,
                           ZN => n8565);
   U9470 : AOI22_X1 port map( A1 => n243, A2 => n5154, B1 => n156, B2 => n5155,
                           ZN => n8564);
   U9471 : NAND3_X1 port map( A1 => n8568, A2 => n8569, A3 => n8570, ZN => 
                           n12419);
   U9472 : AOI221_X1 port map( B1 => n211, B2 => n5159, C1 => n183, C2 => 
                           MEM_IN(29), A => n8571, ZN => n8570);
   U9473 : OAI22_X1 port map( A1 => n11056, A2 => n267, B1 => n5161, B2 => n136
                           , ZN => n8571);
   U9474 : AOI22_X1 port map( A1 => n201, A2 => n5162, B1 => n159, B2 => n5163,
                           ZN => n8569);
   U9475 : AOI22_X1 port map( A1 => n243, A2 => n5164, B1 => n156, B2 => n5165,
                           ZN => n8568);
   U9476 : NAND3_X1 port map( A1 => n8572, A2 => n8573, A3 => n8574, ZN => 
                           n12418);
   U9477 : AOI221_X1 port map( B1 => n211, B2 => n5169, C1 => n183, C2 => 
                           MEM_IN(30), A => n8575, ZN => n8574);
   U9478 : OAI22_X1 port map( A1 => n11055, A2 => n267, B1 => n5171, B2 => n136
                           , ZN => n8575);
   U9479 : AOI22_X1 port map( A1 => n201, A2 => n5172, B1 => n159, B2 => n5173,
                           ZN => n8573);
   U9480 : AOI22_X1 port map( A1 => n243, A2 => n5174, B1 => n156, B2 => n5175,
                           ZN => n8572);
   U9481 : NAND3_X1 port map( A1 => n8576, A2 => n8577, A3 => n8578, ZN => 
                           n12417);
   U9482 : AOI221_X1 port map( B1 => n211, B2 => n5179, C1 => n183, C2 => 
                           MEM_IN(31), A => n8579, ZN => n8578);
   U9483 : OAI22_X1 port map( A1 => n11054, A2 => n267, B1 => n5181, B2 => n136
                           , ZN => n8579);
   U9484 : INV_X1 port map( A => n8585, ZN => n8584);
   U9485 : AOI22_X1 port map( A1 => n201, A2 => n5191, B1 => n159, B2 => n5192,
                           ZN => n8577);
   U9486 : INV_X1 port map( A => n8444, ZN => n8443);
   U9487 : AOI22_X1 port map( A1 => n243, A2 => n5195, B1 => n156, B2 => n5196,
                           ZN => n8576);
   U9488 : AOI22_X1 port map( A1 => n8582, A2 => n8588, B1 => n4841, B2 => n267
                           , ZN => n8583);
   U9489 : INV_X1 port map( A => n8581, ZN => n8588);
   U9490 : NAND3_X1 port map( A1 => n208, A2 => n267, A3 => n7561, ZN => n8581)
                           ;
   U9491 : INV_X1 port map( A => n8580, ZN => n7561);
   U9492 : OAI22_X1 port map( A1 => n8589, A2 => n4786, B1 => n8590, B2 => 
                           n5204, ZN => n8455);
   U9493 : NOR2_X1 port map( A1 => n8580, A2 => n8591, ZN => n8590);
   U9494 : NAND4_X1 port map( A1 => n8447, A2 => n8450, A3 => n7858, A4 => 
                           n7707, ZN => n8580);
   U9495 : NOR4_X1 port map( A1 => n8592, A2 => n8444, A3 => RESET, A4 => n8593
                           , ZN => n8589);
   U9496 : OAI211_X1 port map( C1 => n8594, C2 => n7856, A => n8144, B => n8295
                           , ZN => n8592);
   U9497 : INV_X1 port map( A => n8296, ZN => n8295);
   U9498 : INV_X1 port map( A => n8153, ZN => n8144);
   U9499 : NOR2_X1 port map( A1 => n7707, A2 => n4787, ZN => n8153);
   U9500 : INV_X1 port map( A => n8591, ZN => n8582);
   U9501 : NAND2_X1 port map( A1 => n8595, A2 => n8596, ZN => n8591);
   U9502 : NAND2_X1 port map( A1 => n7708, A2 => n6228, ZN => n7707);
   U9503 : NAND3_X1 port map( A1 => n8597, A2 => n8598, A3 => n8599, ZN => 
                           n12416);
   U9504 : AOI221_X1 port map( B1 => n8600, B2 => n4863, C1 => n184, C2 => 
                           MEM_IN(0), A => n8601, ZN => n8599);
   U9505 : OAI22_X1 port map( A1 => n11053, A2 => n291, B1 => n4867, B2 => n137
                           , ZN => n8601);
   U9506 : AOI22_X1 port map( A1 => n8603, A2 => n4869, B1 => n8604, B2 => 
                           n4871, ZN => n8598);
   U9507 : AOI22_X1 port map( A1 => n8605, A2 => n4873, B1 => n8606, B2 => 
                           n4875, ZN => n8597);
   U9508 : NAND3_X1 port map( A1 => n8607, A2 => n8608, A3 => n8609, ZN => 
                           n12415);
   U9509 : AOI221_X1 port map( B1 => n8600, B2 => n4879, C1 => n184, C2 => 
                           MEM_IN(1), A => n8610, ZN => n8609);
   U9510 : OAI22_X1 port map( A1 => n11052, A2 => n291, B1 => n4881, B2 => n137
                           , ZN => n8610);
   U9511 : AOI22_X1 port map( A1 => n8603, A2 => n4882, B1 => n8604, B2 => 
                           n4883, ZN => n8608);
   U9512 : AOI22_X1 port map( A1 => n8605, A2 => n4884, B1 => n8606, B2 => 
                           n4885, ZN => n8607);
   U9513 : NAND3_X1 port map( A1 => n8611, A2 => n8612, A3 => n8613, ZN => 
                           n12414);
   U9514 : AOI221_X1 port map( B1 => n8600, B2 => n4889, C1 => n184, C2 => 
                           MEM_IN(2), A => n8614, ZN => n8613);
   U9515 : OAI22_X1 port map( A1 => n11051, A2 => n291, B1 => n4891, B2 => n137
                           , ZN => n8614);
   U9516 : AOI22_X1 port map( A1 => n8603, A2 => n4892, B1 => n8604, B2 => 
                           n4893, ZN => n8612);
   U9517 : AOI22_X1 port map( A1 => n8605, A2 => n4894, B1 => n8606, B2 => 
                           n4895, ZN => n8611);
   U9518 : NAND3_X1 port map( A1 => n8615, A2 => n8616, A3 => n8617, ZN => 
                           n12413);
   U9519 : AOI221_X1 port map( B1 => n8600, B2 => n4899, C1 => n184, C2 => 
                           MEM_IN(3), A => n8618, ZN => n8617);
   U9520 : OAI22_X1 port map( A1 => n11050, A2 => n291, B1 => n4901, B2 => n137
                           , ZN => n8618);
   U9521 : AOI22_X1 port map( A1 => n8603, A2 => n4902, B1 => n8604, B2 => 
                           n4903, ZN => n8616);
   U9522 : AOI22_X1 port map( A1 => n8605, A2 => n4904, B1 => n8606, B2 => 
                           n4905, ZN => n8615);
   U9523 : NAND3_X1 port map( A1 => n8619, A2 => n8620, A3 => n8621, ZN => 
                           n12412);
   U9524 : AOI221_X1 port map( B1 => n8600, B2 => n4909, C1 => n184, C2 => 
                           MEM_IN(4), A => n8622, ZN => n8621);
   U9525 : OAI22_X1 port map( A1 => n11049, A2 => n291, B1 => n4911, B2 => n137
                           , ZN => n8622);
   U9526 : AOI22_X1 port map( A1 => n8603, A2 => n4912, B1 => n8604, B2 => 
                           n4913, ZN => n8620);
   U9527 : AOI22_X1 port map( A1 => n8605, A2 => n4914, B1 => n8606, B2 => 
                           n4915, ZN => n8619);
   U9528 : NAND3_X1 port map( A1 => n8623, A2 => n8624, A3 => n8625, ZN => 
                           n12411);
   U9529 : AOI221_X1 port map( B1 => n8600, B2 => n4919, C1 => n184, C2 => 
                           MEM_IN(5), A => n8626, ZN => n8625);
   U9530 : OAI22_X1 port map( A1 => n11048, A2 => n291, B1 => n4921, B2 => n137
                           , ZN => n8626);
   U9531 : AOI22_X1 port map( A1 => n8603, A2 => n4922, B1 => n8604, B2 => 
                           n4923, ZN => n8624);
   U9532 : AOI22_X1 port map( A1 => n8605, A2 => n4924, B1 => n8606, B2 => 
                           n4925, ZN => n8623);
   U9533 : NAND3_X1 port map( A1 => n8627, A2 => n8628, A3 => n8629, ZN => 
                           n12410);
   U9534 : AOI221_X1 port map( B1 => n8600, B2 => n4929, C1 => n184, C2 => 
                           MEM_IN(6), A => n8630, ZN => n8629);
   U9535 : OAI22_X1 port map( A1 => n11047, A2 => n291, B1 => n4931, B2 => n137
                           , ZN => n8630);
   U9536 : AOI22_X1 port map( A1 => n8603, A2 => n4932, B1 => n8604, B2 => 
                           n4933, ZN => n8628);
   U9537 : AOI22_X1 port map( A1 => n8605, A2 => n4934, B1 => n8606, B2 => 
                           n4935, ZN => n8627);
   U9538 : NAND3_X1 port map( A1 => n8631, A2 => n8632, A3 => n8633, ZN => 
                           n12409);
   U9539 : AOI221_X1 port map( B1 => n8600, B2 => n4939, C1 => n184, C2 => 
                           MEM_IN(7), A => n8634, ZN => n8633);
   U9540 : OAI22_X1 port map( A1 => n11046, A2 => n291, B1 => n4941, B2 => n137
                           , ZN => n8634);
   U9541 : AOI22_X1 port map( A1 => n8603, A2 => n4942, B1 => n8604, B2 => 
                           n4943, ZN => n8632);
   U9542 : AOI22_X1 port map( A1 => n8605, A2 => n4944, B1 => n8606, B2 => 
                           n4945, ZN => n8631);
   U9543 : NAND3_X1 port map( A1 => n8635, A2 => n8636, A3 => n8637, ZN => 
                           n12408);
   U9544 : AOI221_X1 port map( B1 => n8600, B2 => n4949, C1 => n184, C2 => 
                           MEM_IN(8), A => n8638, ZN => n8637);
   U9545 : OAI22_X1 port map( A1 => n11045, A2 => n291, B1 => n4951, B2 => n137
                           , ZN => n8638);
   U9546 : AOI22_X1 port map( A1 => n8603, A2 => n4952, B1 => n8604, B2 => 
                           n4953, ZN => n8636);
   U9547 : AOI22_X1 port map( A1 => n8605, A2 => n4954, B1 => n8606, B2 => 
                           n4955, ZN => n8635);
   U9548 : NAND3_X1 port map( A1 => n8639, A2 => n8640, A3 => n8641, ZN => 
                           n12407);
   U9549 : AOI221_X1 port map( B1 => n8600, B2 => n4959, C1 => n184, C2 => 
                           MEM_IN(9), A => n8642, ZN => n8641);
   U9550 : OAI22_X1 port map( A1 => n11044, A2 => n291, B1 => n4961, B2 => n137
                           , ZN => n8642);
   U9551 : AOI22_X1 port map( A1 => n8603, A2 => n4962, B1 => n8604, B2 => 
                           n4963, ZN => n8640);
   U9552 : AOI22_X1 port map( A1 => n8605, A2 => n4964, B1 => n8606, B2 => 
                           n4965, ZN => n8639);
   U9553 : NAND3_X1 port map( A1 => n8643, A2 => n8644, A3 => n8645, ZN => 
                           n12406);
   U9554 : AOI221_X1 port map( B1 => n8600, B2 => n4969, C1 => n184, C2 => 
                           MEM_IN(10), A => n8646, ZN => n8645);
   U9555 : OAI22_X1 port map( A1 => n11043, A2 => n291, B1 => n4971, B2 => n137
                           , ZN => n8646);
   U9556 : AOI22_X1 port map( A1 => n8603, A2 => n4972, B1 => n8604, B2 => 
                           n4973, ZN => n8644);
   U9557 : AOI22_X1 port map( A1 => n8605, A2 => n4974, B1 => n8606, B2 => 
                           n4975, ZN => n8643);
   U9558 : NAND3_X1 port map( A1 => n8647, A2 => n8648, A3 => n8649, ZN => 
                           n12405);
   U9559 : AOI221_X1 port map( B1 => n8600, B2 => n4979, C1 => n184, C2 => 
                           MEM_IN(11), A => n8650, ZN => n8649);
   U9560 : OAI22_X1 port map( A1 => n11042, A2 => n291, B1 => n4981, B2 => n137
                           , ZN => n8650);
   U9561 : AOI22_X1 port map( A1 => n8603, A2 => n4982, B1 => n8604, B2 => 
                           n4983, ZN => n8648);
   U9562 : AOI22_X1 port map( A1 => n8605, A2 => n4984, B1 => n8606, B2 => 
                           n4985, ZN => n8647);
   U9563 : NAND3_X1 port map( A1 => n8651, A2 => n8652, A3 => n8653, ZN => 
                           n12404);
   U9564 : AOI221_X1 port map( B1 => n8600, B2 => n4989, C1 => n184, C2 => 
                           MEM_IN(12), A => n8654, ZN => n8653);
   U9565 : OAI22_X1 port map( A1 => n11041, A2 => n291, B1 => n4991, B2 => n137
                           , ZN => n8654);
   U9566 : AOI22_X1 port map( A1 => n8603, A2 => n4992, B1 => n8604, B2 => 
                           n4993, ZN => n8652);
   U9567 : AOI22_X1 port map( A1 => n8605, A2 => n4994, B1 => n8606, B2 => 
                           n4995, ZN => n8651);
   U9568 : NAND3_X1 port map( A1 => n8655, A2 => n8656, A3 => n8657, ZN => 
                           n12403);
   U9569 : AOI221_X1 port map( B1 => n8600, B2 => n4999, C1 => n184, C2 => 
                           MEM_IN(13), A => n8658, ZN => n8657);
   U9570 : OAI22_X1 port map( A1 => n11040, A2 => n291, B1 => n5001, B2 => n137
                           , ZN => n8658);
   U9571 : AOI22_X1 port map( A1 => n8603, A2 => n5002, B1 => n8604, B2 => 
                           n5003, ZN => n8656);
   U9572 : AOI22_X1 port map( A1 => n8605, A2 => n5004, B1 => n8606, B2 => 
                           n5005, ZN => n8655);
   U9573 : NAND3_X1 port map( A1 => n8659, A2 => n8660, A3 => n8661, ZN => 
                           n12402);
   U9574 : AOI221_X1 port map( B1 => n8600, B2 => n5009, C1 => n184, C2 => 
                           MEM_IN(14), A => n8662, ZN => n8661);
   U9575 : OAI22_X1 port map( A1 => n11039, A2 => n291, B1 => n5011, B2 => n137
                           , ZN => n8662);
   U9576 : AOI22_X1 port map( A1 => n8603, A2 => n5012, B1 => n8604, B2 => 
                           n5013, ZN => n8660);
   U9577 : AOI22_X1 port map( A1 => n8605, A2 => n5014, B1 => n8606, B2 => 
                           n5015, ZN => n8659);
   U9578 : NAND3_X1 port map( A1 => n8663, A2 => n8664, A3 => n8665, ZN => 
                           n12401);
   U9579 : AOI221_X1 port map( B1 => n8600, B2 => n5019, C1 => n184, C2 => 
                           MEM_IN(15), A => n8666, ZN => n8665);
   U9580 : OAI22_X1 port map( A1 => n11038, A2 => n291, B1 => n5021, B2 => n137
                           , ZN => n8666);
   U9581 : AOI22_X1 port map( A1 => n8603, A2 => n5022, B1 => n8604, B2 => 
                           n5023, ZN => n8664);
   U9582 : AOI22_X1 port map( A1 => n8605, A2 => n5024, B1 => n8606, B2 => 
                           n5025, ZN => n8663);
   U9583 : NAND3_X1 port map( A1 => n8667, A2 => n8668, A3 => n8669, ZN => 
                           n12400);
   U9584 : AOI221_X1 port map( B1 => n8600, B2 => n5029, C1 => n184, C2 => 
                           MEM_IN(16), A => n8670, ZN => n8669);
   U9585 : OAI22_X1 port map( A1 => n11037, A2 => n291, B1 => n5031, B2 => n137
                           , ZN => n8670);
   U9586 : AOI22_X1 port map( A1 => n8603, A2 => n5032, B1 => n8604, B2 => 
                           n5033, ZN => n8668);
   U9587 : AOI22_X1 port map( A1 => n8605, A2 => n5034, B1 => n8606, B2 => 
                           n5035, ZN => n8667);
   U9588 : NAND3_X1 port map( A1 => n8671, A2 => n8672, A3 => n8673, ZN => 
                           n12399);
   U9589 : AOI221_X1 port map( B1 => n8600, B2 => n5039, C1 => n184, C2 => 
                           MEM_IN(17), A => n8674, ZN => n8673);
   U9590 : OAI22_X1 port map( A1 => n11036, A2 => n291, B1 => n5041, B2 => n137
                           , ZN => n8674);
   U9591 : AOI22_X1 port map( A1 => n8603, A2 => n5042, B1 => n8604, B2 => 
                           n5043, ZN => n8672);
   U9592 : AOI22_X1 port map( A1 => n8605, A2 => n5044, B1 => n8606, B2 => 
                           n5045, ZN => n8671);
   U9593 : NAND3_X1 port map( A1 => n8675, A2 => n8676, A3 => n8677, ZN => 
                           n12398);
   U9594 : AOI221_X1 port map( B1 => n8600, B2 => n5049, C1 => n184, C2 => 
                           MEM_IN(18), A => n8678, ZN => n8677);
   U9595 : OAI22_X1 port map( A1 => n11035, A2 => n291, B1 => n5051, B2 => n137
                           , ZN => n8678);
   U9596 : AOI22_X1 port map( A1 => n8603, A2 => n5052, B1 => n8604, B2 => 
                           n5053, ZN => n8676);
   U9597 : AOI22_X1 port map( A1 => n8605, A2 => n5054, B1 => n8606, B2 => 
                           n5055, ZN => n8675);
   U9598 : NAND3_X1 port map( A1 => n8679, A2 => n8680, A3 => n8681, ZN => 
                           n12397);
   U9599 : AOI221_X1 port map( B1 => n8600, B2 => n5059, C1 => n184, C2 => 
                           MEM_IN(19), A => n8682, ZN => n8681);
   U9600 : OAI22_X1 port map( A1 => n11034, A2 => n291, B1 => n5061, B2 => n137
                           , ZN => n8682);
   U9601 : AOI22_X1 port map( A1 => n8603, A2 => n5062, B1 => n8604, B2 => 
                           n5063, ZN => n8680);
   U9602 : AOI22_X1 port map( A1 => n8605, A2 => n5064, B1 => n8606, B2 => 
                           n5065, ZN => n8679);
   U9603 : NAND3_X1 port map( A1 => n8683, A2 => n8684, A3 => n8685, ZN => 
                           n12396);
   U9604 : AOI221_X1 port map( B1 => n8600, B2 => n5069, C1 => n184, C2 => 
                           MEM_IN(20), A => n8686, ZN => n8685);
   U9605 : OAI22_X1 port map( A1 => n11033, A2 => n291, B1 => n5071, B2 => n137
                           , ZN => n8686);
   U9606 : AOI22_X1 port map( A1 => n8603, A2 => n5072, B1 => n8604, B2 => 
                           n5073, ZN => n8684);
   U9607 : AOI22_X1 port map( A1 => n8605, A2 => n5074, B1 => n8606, B2 => 
                           n5075, ZN => n8683);
   U9608 : NAND3_X1 port map( A1 => n8687, A2 => n8688, A3 => n8689, ZN => 
                           n12395);
   U9609 : AOI221_X1 port map( B1 => n8600, B2 => n5079, C1 => n184, C2 => 
                           MEM_IN(21), A => n8690, ZN => n8689);
   U9610 : OAI22_X1 port map( A1 => n11032, A2 => n291, B1 => n5081, B2 => n137
                           , ZN => n8690);
   U9611 : AOI22_X1 port map( A1 => n8603, A2 => n5082, B1 => n8604, B2 => 
                           n5083, ZN => n8688);
   U9612 : AOI22_X1 port map( A1 => n8605, A2 => n5084, B1 => n8606, B2 => 
                           n5085, ZN => n8687);
   U9613 : NAND3_X1 port map( A1 => n8691, A2 => n8692, A3 => n8693, ZN => 
                           n12394);
   U9614 : AOI221_X1 port map( B1 => n8600, B2 => n5089, C1 => n184, C2 => 
                           MEM_IN(22), A => n8694, ZN => n8693);
   U9615 : OAI22_X1 port map( A1 => n11031, A2 => n291, B1 => n5091, B2 => n137
                           , ZN => n8694);
   U9616 : AOI22_X1 port map( A1 => n8603, A2 => n5092, B1 => n8604, B2 => 
                           n5093, ZN => n8692);
   U9617 : AOI22_X1 port map( A1 => n8605, A2 => n5094, B1 => n8606, B2 => 
                           n5095, ZN => n8691);
   U9618 : NAND3_X1 port map( A1 => n8695, A2 => n8696, A3 => n8697, ZN => 
                           n12393);
   U9619 : AOI221_X1 port map( B1 => n8600, B2 => n5099, C1 => n184, C2 => 
                           MEM_IN(23), A => n8698, ZN => n8697);
   U9620 : OAI22_X1 port map( A1 => n11030, A2 => n291, B1 => n5101, B2 => n137
                           , ZN => n8698);
   U9621 : AOI22_X1 port map( A1 => n8603, A2 => n5102, B1 => n8604, B2 => 
                           n5103, ZN => n8696);
   U9622 : AOI22_X1 port map( A1 => n8605, A2 => n5104, B1 => n8606, B2 => 
                           n5105, ZN => n8695);
   U9623 : NAND3_X1 port map( A1 => n8699, A2 => n8700, A3 => n8701, ZN => 
                           n12392);
   U9624 : AOI221_X1 port map( B1 => n8600, B2 => n5109, C1 => n184, C2 => 
                           MEM_IN(24), A => n8702, ZN => n8701);
   U9625 : OAI22_X1 port map( A1 => n11029, A2 => n291, B1 => n5111, B2 => n137
                           , ZN => n8702);
   U9626 : AOI22_X1 port map( A1 => n8603, A2 => n5112, B1 => n8604, B2 => 
                           n5113, ZN => n8700);
   U9627 : AOI22_X1 port map( A1 => n8605, A2 => n5114, B1 => n8606, B2 => 
                           n5115, ZN => n8699);
   U9628 : NAND3_X1 port map( A1 => n8703, A2 => n8704, A3 => n8705, ZN => 
                           n12391);
   U9629 : AOI221_X1 port map( B1 => n8600, B2 => n5119, C1 => n184, C2 => 
                           MEM_IN(25), A => n8706, ZN => n8705);
   U9630 : OAI22_X1 port map( A1 => n11028, A2 => n291, B1 => n5121, B2 => n137
                           , ZN => n8706);
   U9631 : AOI22_X1 port map( A1 => n8603, A2 => n5122, B1 => n8604, B2 => 
                           n5123, ZN => n8704);
   U9632 : AOI22_X1 port map( A1 => n8605, A2 => n5124, B1 => n8606, B2 => 
                           n5125, ZN => n8703);
   U9633 : NAND3_X1 port map( A1 => n8707, A2 => n8708, A3 => n8709, ZN => 
                           n12390);
   U9634 : AOI221_X1 port map( B1 => n8600, B2 => n5129, C1 => n184, C2 => 
                           MEM_IN(26), A => n8710, ZN => n8709);
   U9635 : OAI22_X1 port map( A1 => n11027, A2 => n291, B1 => n5131, B2 => n137
                           , ZN => n8710);
   U9636 : AOI22_X1 port map( A1 => n8603, A2 => n5132, B1 => n8604, B2 => 
                           n5133, ZN => n8708);
   U9637 : AOI22_X1 port map( A1 => n8605, A2 => n5134, B1 => n8606, B2 => 
                           n5135, ZN => n8707);
   U9638 : NAND3_X1 port map( A1 => n8711, A2 => n8712, A3 => n8713, ZN => 
                           n12389);
   U9639 : AOI221_X1 port map( B1 => n8600, B2 => n5139, C1 => n184, C2 => 
                           MEM_IN(27), A => n8714, ZN => n8713);
   U9640 : OAI22_X1 port map( A1 => n11026, A2 => n291, B1 => n5141, B2 => n137
                           , ZN => n8714);
   U9641 : AOI22_X1 port map( A1 => n8603, A2 => n5142, B1 => n8604, B2 => 
                           n5143, ZN => n8712);
   U9642 : AOI22_X1 port map( A1 => n8605, A2 => n5144, B1 => n8606, B2 => 
                           n5145, ZN => n8711);
   U9643 : NAND3_X1 port map( A1 => n8715, A2 => n8716, A3 => n8717, ZN => 
                           n12388);
   U9644 : AOI221_X1 port map( B1 => n8600, B2 => n5149, C1 => n184, C2 => 
                           MEM_IN(28), A => n8718, ZN => n8717);
   U9645 : OAI22_X1 port map( A1 => n11025, A2 => n291, B1 => n5151, B2 => n137
                           , ZN => n8718);
   U9646 : AOI22_X1 port map( A1 => n8603, A2 => n5152, B1 => n8604, B2 => 
                           n5153, ZN => n8716);
   U9647 : AOI22_X1 port map( A1 => n8605, A2 => n5154, B1 => n8606, B2 => 
                           n5155, ZN => n8715);
   U9648 : NAND3_X1 port map( A1 => n8719, A2 => n8720, A3 => n8721, ZN => 
                           n12387);
   U9649 : AOI221_X1 port map( B1 => n8600, B2 => n5159, C1 => n184, C2 => 
                           MEM_IN(29), A => n8722, ZN => n8721);
   U9650 : OAI22_X1 port map( A1 => n11024, A2 => n291, B1 => n5161, B2 => n137
                           , ZN => n8722);
   U9651 : AOI22_X1 port map( A1 => n8603, A2 => n5162, B1 => n8604, B2 => 
                           n5163, ZN => n8720);
   U9652 : AOI22_X1 port map( A1 => n8605, A2 => n5164, B1 => n8606, B2 => 
                           n5165, ZN => n8719);
   U9653 : NAND3_X1 port map( A1 => n8723, A2 => n8724, A3 => n8725, ZN => 
                           n12386);
   U9654 : AOI221_X1 port map( B1 => n8600, B2 => n5169, C1 => n184, C2 => 
                           MEM_IN(30), A => n8726, ZN => n8725);
   U9655 : OAI22_X1 port map( A1 => n11023, A2 => n291, B1 => n5171, B2 => n137
                           , ZN => n8726);
   U9656 : AOI22_X1 port map( A1 => n8603, A2 => n5172, B1 => n8604, B2 => 
                           n5173, ZN => n8724);
   U9657 : AOI22_X1 port map( A1 => n8605, A2 => n5174, B1 => n8606, B2 => 
                           n5175, ZN => n8723);
   U9658 : NAND3_X1 port map( A1 => n8727, A2 => n8728, A3 => n8729, ZN => 
                           n12385);
   U9659 : AOI221_X1 port map( B1 => n8600, B2 => n5179, C1 => n184, C2 => 
                           MEM_IN(31), A => n8730, ZN => n8729);
   U9660 : OAI22_X1 port map( A1 => n11022, A2 => n291, B1 => n5181, B2 => n137
                           , ZN => n8730);
   U9661 : INV_X1 port map( A => n8734, ZN => n8733);
   U9662 : NAND2_X1 port map( A1 => n5206, A2 => n8587, ZN => n8585);
   U9663 : NAND3_X1 port map( A1 => n5206, A2 => n7858, A3 => n8299, ZN => 
                           n8587);
   U9664 : AOI22_X1 port map( A1 => n8603, A2 => n5191, B1 => n8604, B2 => 
                           n5192, ZN => n8728);
   U9665 : AOI22_X1 port map( A1 => n8605, A2 => n5195, B1 => n8606, B2 => 
                           n5196, ZN => n8727);
   U9666 : OAI22_X1 port map( A1 => n8734, A2 => n8732, B1 => n208, B2 => n290,
                           ZN => n8736);
   U9667 : NAND3_X1 port map( A1 => n208, A2 => n291, A3 => n7706, ZN => n8732)
                           ;
   U9668 : INV_X1 port map( A => n8731, ZN => n7706);
   U9669 : OAI22_X1 port map( A1 => n4786, A2 => n8738, B1 => n8739, B2 => 
                           n5204, ZN => n8602);
   U9670 : NOR2_X1 port map( A1 => n8731, A2 => n8734, ZN => n8739);
   U9671 : NAND3_X1 port map( A1 => n8447, A2 => n7858, A3 => n8740, ZN => 
                           n8731);
   U9672 : NOR3_X1 port map( A1 => n8741, A2 => RESET, A3 => n8296, ZN => n8738
                           );
   U9673 : OAI22_X1 port map( A1 => n8447, A2 => n4787, B1 => n6374, B2 => 
                           n7856, ZN => n8741);
   U9674 : NAND3_X1 port map( A1 => n6378, A2 => n8742, A3 => n7560, ZN => 
                           n7856);
   U9675 : INV_X1 port map( A => n8743, ZN => n6378);
   U9676 : NAND2_X1 port map( A1 => n8744, A2 => n8745, ZN => n8734);
   U9677 : NOR2_X1 port map( A1 => n7858, A2 => n4787, ZN => n8296);
   U9678 : NAND2_X1 port map( A1 => n7708, A2 => n6381, ZN => n7858);
   U9679 : NAND3_X1 port map( A1 => n8746, A2 => n8747, A3 => n8748, ZN => 
                           n12384);
   U9680 : AOI221_X1 port map( B1 => n8749, B2 => n4863, C1 => n185, C2 => 
                           MEM_IN(0), A => n8750, ZN => n8748);
   U9681 : OAI22_X1 port map( A1 => n11021, A2 => n277, B1 => n4867, B2 => n134
                           , ZN => n8750);
   U9682 : AOI22_X1 port map( A1 => n8752, A2 => n4869, B1 => n8753, B2 => 
                           n4871, ZN => n8747);
   U9683 : AOI22_X1 port map( A1 => n8754, A2 => n4873, B1 => n8755, B2 => 
                           n4875, ZN => n8746);
   U9684 : NAND3_X1 port map( A1 => n8756, A2 => n8757, A3 => n8758, ZN => 
                           n12383);
   U9685 : AOI221_X1 port map( B1 => n8749, B2 => n4879, C1 => n185, C2 => 
                           MEM_IN(1), A => n8759, ZN => n8758);
   U9686 : OAI22_X1 port map( A1 => n11020, A2 => n277, B1 => n4881, B2 => n134
                           , ZN => n8759);
   U9687 : AOI22_X1 port map( A1 => n8752, A2 => n4882, B1 => n8753, B2 => 
                           n4883, ZN => n8757);
   U9688 : AOI22_X1 port map( A1 => n8754, A2 => n4884, B1 => n8755, B2 => 
                           n4885, ZN => n8756);
   U9689 : NAND3_X1 port map( A1 => n8760, A2 => n8761, A3 => n8762, ZN => 
                           n12382);
   U9690 : AOI221_X1 port map( B1 => n8749, B2 => n4889, C1 => n185, C2 => 
                           MEM_IN(2), A => n8763, ZN => n8762);
   U9691 : OAI22_X1 port map( A1 => n11019, A2 => n277, B1 => n4891, B2 => n134
                           , ZN => n8763);
   U9692 : AOI22_X1 port map( A1 => n8752, A2 => n4892, B1 => n8753, B2 => 
                           n4893, ZN => n8761);
   U9693 : AOI22_X1 port map( A1 => n8754, A2 => n4894, B1 => n8755, B2 => 
                           n4895, ZN => n8760);
   U9694 : NAND3_X1 port map( A1 => n8764, A2 => n8765, A3 => n8766, ZN => 
                           n12381);
   U9695 : AOI221_X1 port map( B1 => n8749, B2 => n4899, C1 => n185, C2 => 
                           MEM_IN(3), A => n8767, ZN => n8766);
   U9696 : OAI22_X1 port map( A1 => n11018, A2 => n277, B1 => n4901, B2 => n134
                           , ZN => n8767);
   U9697 : AOI22_X1 port map( A1 => n8752, A2 => n4902, B1 => n8753, B2 => 
                           n4903, ZN => n8765);
   U9698 : AOI22_X1 port map( A1 => n8754, A2 => n4904, B1 => n8755, B2 => 
                           n4905, ZN => n8764);
   U9699 : NAND3_X1 port map( A1 => n8768, A2 => n8769, A3 => n8770, ZN => 
                           n12380);
   U9700 : AOI221_X1 port map( B1 => n8749, B2 => n4909, C1 => n185, C2 => 
                           MEM_IN(4), A => n8771, ZN => n8770);
   U9701 : OAI22_X1 port map( A1 => n11017, A2 => n277, B1 => n4911, B2 => n134
                           , ZN => n8771);
   U9702 : AOI22_X1 port map( A1 => n8752, A2 => n4912, B1 => n8753, B2 => 
                           n4913, ZN => n8769);
   U9703 : AOI22_X1 port map( A1 => n8754, A2 => n4914, B1 => n8755, B2 => 
                           n4915, ZN => n8768);
   U9704 : NAND3_X1 port map( A1 => n8772, A2 => n8773, A3 => n8774, ZN => 
                           n12379);
   U9705 : AOI221_X1 port map( B1 => n8749, B2 => n4919, C1 => n185, C2 => 
                           MEM_IN(5), A => n8775, ZN => n8774);
   U9706 : OAI22_X1 port map( A1 => n11016, A2 => n277, B1 => n4921, B2 => n134
                           , ZN => n8775);
   U9707 : AOI22_X1 port map( A1 => n8752, A2 => n4922, B1 => n8753, B2 => 
                           n4923, ZN => n8773);
   U9708 : AOI22_X1 port map( A1 => n8754, A2 => n4924, B1 => n8755, B2 => 
                           n4925, ZN => n8772);
   U9709 : NAND3_X1 port map( A1 => n8776, A2 => n8777, A3 => n8778, ZN => 
                           n12378);
   U9710 : AOI221_X1 port map( B1 => n8749, B2 => n4929, C1 => n185, C2 => 
                           MEM_IN(6), A => n8779, ZN => n8778);
   U9711 : OAI22_X1 port map( A1 => n11015, A2 => n277, B1 => n4931, B2 => n134
                           , ZN => n8779);
   U9712 : AOI22_X1 port map( A1 => n8752, A2 => n4932, B1 => n8753, B2 => 
                           n4933, ZN => n8777);
   U9713 : AOI22_X1 port map( A1 => n8754, A2 => n4934, B1 => n8755, B2 => 
                           n4935, ZN => n8776);
   U9714 : NAND3_X1 port map( A1 => n8780, A2 => n8781, A3 => n8782, ZN => 
                           n12377);
   U9715 : AOI221_X1 port map( B1 => n8749, B2 => n4939, C1 => n185, C2 => 
                           MEM_IN(7), A => n8783, ZN => n8782);
   U9716 : OAI22_X1 port map( A1 => n11014, A2 => n277, B1 => n4941, B2 => n134
                           , ZN => n8783);
   U9717 : AOI22_X1 port map( A1 => n8752, A2 => n4942, B1 => n8753, B2 => 
                           n4943, ZN => n8781);
   U9718 : AOI22_X1 port map( A1 => n8754, A2 => n4944, B1 => n8755, B2 => 
                           n4945, ZN => n8780);
   U9719 : NAND3_X1 port map( A1 => n8784, A2 => n8785, A3 => n8786, ZN => 
                           n12376);
   U9720 : AOI221_X1 port map( B1 => n8749, B2 => n4949, C1 => n185, C2 => 
                           MEM_IN(8), A => n8787, ZN => n8786);
   U9721 : OAI22_X1 port map( A1 => n11013, A2 => n277, B1 => n4951, B2 => n134
                           , ZN => n8787);
   U9722 : AOI22_X1 port map( A1 => n8752, A2 => n4952, B1 => n8753, B2 => 
                           n4953, ZN => n8785);
   U9723 : AOI22_X1 port map( A1 => n8754, A2 => n4954, B1 => n8755, B2 => 
                           n4955, ZN => n8784);
   U9724 : NAND3_X1 port map( A1 => n8788, A2 => n8789, A3 => n8790, ZN => 
                           n12375);
   U9725 : AOI221_X1 port map( B1 => n8749, B2 => n4959, C1 => n185, C2 => 
                           MEM_IN(9), A => n8791, ZN => n8790);
   U9726 : OAI22_X1 port map( A1 => n11012, A2 => n277, B1 => n4961, B2 => n134
                           , ZN => n8791);
   U9727 : AOI22_X1 port map( A1 => n8752, A2 => n4962, B1 => n8753, B2 => 
                           n4963, ZN => n8789);
   U9728 : AOI22_X1 port map( A1 => n8754, A2 => n4964, B1 => n8755, B2 => 
                           n4965, ZN => n8788);
   U9729 : NAND3_X1 port map( A1 => n8792, A2 => n8793, A3 => n8794, ZN => 
                           n12374);
   U9730 : AOI221_X1 port map( B1 => n8749, B2 => n4969, C1 => n185, C2 => 
                           MEM_IN(10), A => n8795, ZN => n8794);
   U9731 : OAI22_X1 port map( A1 => n11011, A2 => n277, B1 => n4971, B2 => n134
                           , ZN => n8795);
   U9732 : AOI22_X1 port map( A1 => n8752, A2 => n4972, B1 => n8753, B2 => 
                           n4973, ZN => n8793);
   U9733 : AOI22_X1 port map( A1 => n8754, A2 => n4974, B1 => n8755, B2 => 
                           n4975, ZN => n8792);
   U9734 : NAND3_X1 port map( A1 => n8796, A2 => n8797, A3 => n8798, ZN => 
                           n12373);
   U9735 : AOI221_X1 port map( B1 => n8749, B2 => n4979, C1 => n185, C2 => 
                           MEM_IN(11), A => n8799, ZN => n8798);
   U9736 : OAI22_X1 port map( A1 => n11010, A2 => n277, B1 => n4981, B2 => n134
                           , ZN => n8799);
   U9737 : AOI22_X1 port map( A1 => n8752, A2 => n4982, B1 => n8753, B2 => 
                           n4983, ZN => n8797);
   U9738 : AOI22_X1 port map( A1 => n8754, A2 => n4984, B1 => n8755, B2 => 
                           n4985, ZN => n8796);
   U9739 : NAND3_X1 port map( A1 => n8800, A2 => n8801, A3 => n8802, ZN => 
                           n12372);
   U9740 : AOI221_X1 port map( B1 => n8749, B2 => n4989, C1 => n185, C2 => 
                           MEM_IN(12), A => n8803, ZN => n8802);
   U9741 : OAI22_X1 port map( A1 => n11009, A2 => n277, B1 => n4991, B2 => n134
                           , ZN => n8803);
   U9742 : AOI22_X1 port map( A1 => n8752, A2 => n4992, B1 => n8753, B2 => 
                           n4993, ZN => n8801);
   U9743 : AOI22_X1 port map( A1 => n8754, A2 => n4994, B1 => n8755, B2 => 
                           n4995, ZN => n8800);
   U9744 : NAND3_X1 port map( A1 => n8804, A2 => n8805, A3 => n8806, ZN => 
                           n12371);
   U9745 : AOI221_X1 port map( B1 => n8749, B2 => n4999, C1 => n185, C2 => 
                           MEM_IN(13), A => n8807, ZN => n8806);
   U9746 : OAI22_X1 port map( A1 => n11008, A2 => n277, B1 => n5001, B2 => n134
                           , ZN => n8807);
   U9747 : AOI22_X1 port map( A1 => n8752, A2 => n5002, B1 => n8753, B2 => 
                           n5003, ZN => n8805);
   U9748 : AOI22_X1 port map( A1 => n8754, A2 => n5004, B1 => n8755, B2 => 
                           n5005, ZN => n8804);
   U9749 : NAND3_X1 port map( A1 => n8808, A2 => n8809, A3 => n8810, ZN => 
                           n12370);
   U9750 : AOI221_X1 port map( B1 => n8749, B2 => n5009, C1 => n185, C2 => 
                           MEM_IN(14), A => n8811, ZN => n8810);
   U9751 : OAI22_X1 port map( A1 => n11007, A2 => n277, B1 => n5011, B2 => n134
                           , ZN => n8811);
   U9752 : AOI22_X1 port map( A1 => n8752, A2 => n5012, B1 => n8753, B2 => 
                           n5013, ZN => n8809);
   U9753 : AOI22_X1 port map( A1 => n8754, A2 => n5014, B1 => n8755, B2 => 
                           n5015, ZN => n8808);
   U9754 : NAND3_X1 port map( A1 => n8812, A2 => n8813, A3 => n8814, ZN => 
                           n12369);
   U9755 : AOI221_X1 port map( B1 => n8749, B2 => n5019, C1 => n185, C2 => 
                           MEM_IN(15), A => n8815, ZN => n8814);
   U9756 : OAI22_X1 port map( A1 => n11006, A2 => n277, B1 => n5021, B2 => n134
                           , ZN => n8815);
   U9757 : AOI22_X1 port map( A1 => n8752, A2 => n5022, B1 => n8753, B2 => 
                           n5023, ZN => n8813);
   U9758 : AOI22_X1 port map( A1 => n8754, A2 => n5024, B1 => n8755, B2 => 
                           n5025, ZN => n8812);
   U9759 : NAND3_X1 port map( A1 => n8816, A2 => n8817, A3 => n8818, ZN => 
                           n12368);
   U9760 : AOI221_X1 port map( B1 => n8749, B2 => n5029, C1 => n185, C2 => 
                           MEM_IN(16), A => n8819, ZN => n8818);
   U9761 : OAI22_X1 port map( A1 => n11005, A2 => n277, B1 => n5031, B2 => n134
                           , ZN => n8819);
   U9762 : AOI22_X1 port map( A1 => n8752, A2 => n5032, B1 => n8753, B2 => 
                           n5033, ZN => n8817);
   U9763 : AOI22_X1 port map( A1 => n8754, A2 => n5034, B1 => n8755, B2 => 
                           n5035, ZN => n8816);
   U9764 : NAND3_X1 port map( A1 => n8820, A2 => n8821, A3 => n8822, ZN => 
                           n12367);
   U9765 : AOI221_X1 port map( B1 => n8749, B2 => n5039, C1 => n185, C2 => 
                           MEM_IN(17), A => n8823, ZN => n8822);
   U9766 : OAI22_X1 port map( A1 => n11004, A2 => n277, B1 => n5041, B2 => n134
                           , ZN => n8823);
   U9767 : AOI22_X1 port map( A1 => n8752, A2 => n5042, B1 => n8753, B2 => 
                           n5043, ZN => n8821);
   U9768 : AOI22_X1 port map( A1 => n8754, A2 => n5044, B1 => n8755, B2 => 
                           n5045, ZN => n8820);
   U9769 : NAND3_X1 port map( A1 => n8824, A2 => n8825, A3 => n8826, ZN => 
                           n12366);
   U9770 : AOI221_X1 port map( B1 => n8749, B2 => n5049, C1 => n185, C2 => 
                           MEM_IN(18), A => n8827, ZN => n8826);
   U9771 : OAI22_X1 port map( A1 => n11003, A2 => n277, B1 => n5051, B2 => n134
                           , ZN => n8827);
   U9772 : AOI22_X1 port map( A1 => n8752, A2 => n5052, B1 => n8753, B2 => 
                           n5053, ZN => n8825);
   U9773 : AOI22_X1 port map( A1 => n8754, A2 => n5054, B1 => n8755, B2 => 
                           n5055, ZN => n8824);
   U9774 : NAND3_X1 port map( A1 => n8828, A2 => n8829, A3 => n8830, ZN => 
                           n12365);
   U9775 : AOI221_X1 port map( B1 => n8749, B2 => n5059, C1 => n185, C2 => 
                           MEM_IN(19), A => n8831, ZN => n8830);
   U9776 : OAI22_X1 port map( A1 => n11002, A2 => n277, B1 => n5061, B2 => n134
                           , ZN => n8831);
   U9777 : AOI22_X1 port map( A1 => n8752, A2 => n5062, B1 => n8753, B2 => 
                           n5063, ZN => n8829);
   U9778 : AOI22_X1 port map( A1 => n8754, A2 => n5064, B1 => n8755, B2 => 
                           n5065, ZN => n8828);
   U9779 : NAND3_X1 port map( A1 => n8832, A2 => n8833, A3 => n8834, ZN => 
                           n12364);
   U9780 : AOI221_X1 port map( B1 => n8749, B2 => n5069, C1 => n185, C2 => 
                           MEM_IN(20), A => n8835, ZN => n8834);
   U9781 : OAI22_X1 port map( A1 => n11001, A2 => n277, B1 => n5071, B2 => n134
                           , ZN => n8835);
   U9782 : AOI22_X1 port map( A1 => n8752, A2 => n5072, B1 => n8753, B2 => 
                           n5073, ZN => n8833);
   U9783 : AOI22_X1 port map( A1 => n8754, A2 => n5074, B1 => n8755, B2 => 
                           n5075, ZN => n8832);
   U9784 : NAND3_X1 port map( A1 => n8836, A2 => n8837, A3 => n8838, ZN => 
                           n12363);
   U9785 : AOI221_X1 port map( B1 => n8749, B2 => n5079, C1 => n185, C2 => 
                           MEM_IN(21), A => n8839, ZN => n8838);
   U9786 : OAI22_X1 port map( A1 => n11000, A2 => n277, B1 => n5081, B2 => n134
                           , ZN => n8839);
   U9787 : AOI22_X1 port map( A1 => n8752, A2 => n5082, B1 => n8753, B2 => 
                           n5083, ZN => n8837);
   U9788 : AOI22_X1 port map( A1 => n8754, A2 => n5084, B1 => n8755, B2 => 
                           n5085, ZN => n8836);
   U9789 : NAND3_X1 port map( A1 => n8840, A2 => n8841, A3 => n8842, ZN => 
                           n12362);
   U9790 : AOI221_X1 port map( B1 => n8749, B2 => n5089, C1 => n185, C2 => 
                           MEM_IN(22), A => n8843, ZN => n8842);
   U9791 : OAI22_X1 port map( A1 => n10999, A2 => n277, B1 => n5091, B2 => n134
                           , ZN => n8843);
   U9792 : AOI22_X1 port map( A1 => n8752, A2 => n5092, B1 => n8753, B2 => 
                           n5093, ZN => n8841);
   U9793 : AOI22_X1 port map( A1 => n8754, A2 => n5094, B1 => n8755, B2 => 
                           n5095, ZN => n8840);
   U9794 : NAND3_X1 port map( A1 => n8844, A2 => n8845, A3 => n8846, ZN => 
                           n12361);
   U9795 : AOI221_X1 port map( B1 => n8749, B2 => n5099, C1 => n185, C2 => 
                           MEM_IN(23), A => n8847, ZN => n8846);
   U9796 : OAI22_X1 port map( A1 => n10998, A2 => n277, B1 => n5101, B2 => n134
                           , ZN => n8847);
   U9797 : AOI22_X1 port map( A1 => n8752, A2 => n5102, B1 => n8753, B2 => 
                           n5103, ZN => n8845);
   U9798 : AOI22_X1 port map( A1 => n8754, A2 => n5104, B1 => n8755, B2 => 
                           n5105, ZN => n8844);
   U9799 : NAND3_X1 port map( A1 => n8848, A2 => n8849, A3 => n8850, ZN => 
                           n12360);
   U9800 : AOI221_X1 port map( B1 => n8749, B2 => n5109, C1 => n185, C2 => 
                           MEM_IN(24), A => n8851, ZN => n8850);
   U9801 : OAI22_X1 port map( A1 => n10997, A2 => n277, B1 => n5111, B2 => n134
                           , ZN => n8851);
   U9802 : AOI22_X1 port map( A1 => n8752, A2 => n5112, B1 => n8753, B2 => 
                           n5113, ZN => n8849);
   U9803 : AOI22_X1 port map( A1 => n8754, A2 => n5114, B1 => n8755, B2 => 
                           n5115, ZN => n8848);
   U9804 : NAND3_X1 port map( A1 => n8852, A2 => n8853, A3 => n8854, ZN => 
                           n12359);
   U9805 : AOI221_X1 port map( B1 => n8749, B2 => n5119, C1 => n185, C2 => 
                           MEM_IN(25), A => n8855, ZN => n8854);
   U9806 : OAI22_X1 port map( A1 => n10996, A2 => n277, B1 => n5121, B2 => n134
                           , ZN => n8855);
   U9807 : AOI22_X1 port map( A1 => n8752, A2 => n5122, B1 => n8753, B2 => 
                           n5123, ZN => n8853);
   U9808 : AOI22_X1 port map( A1 => n8754, A2 => n5124, B1 => n8755, B2 => 
                           n5125, ZN => n8852);
   U9809 : NAND3_X1 port map( A1 => n8856, A2 => n8857, A3 => n8858, ZN => 
                           n12358);
   U9810 : AOI221_X1 port map( B1 => n8749, B2 => n5129, C1 => n185, C2 => 
                           MEM_IN(26), A => n8859, ZN => n8858);
   U9811 : OAI22_X1 port map( A1 => n10995, A2 => n277, B1 => n5131, B2 => n134
                           , ZN => n8859);
   U9812 : AOI22_X1 port map( A1 => n8752, A2 => n5132, B1 => n8753, B2 => 
                           n5133, ZN => n8857);
   U9813 : AOI22_X1 port map( A1 => n8754, A2 => n5134, B1 => n8755, B2 => 
                           n5135, ZN => n8856);
   U9814 : NAND3_X1 port map( A1 => n8860, A2 => n8861, A3 => n8862, ZN => 
                           n12357);
   U9815 : AOI221_X1 port map( B1 => n8749, B2 => n5139, C1 => n185, C2 => 
                           MEM_IN(27), A => n8863, ZN => n8862);
   U9816 : OAI22_X1 port map( A1 => n10994, A2 => n277, B1 => n5141, B2 => n134
                           , ZN => n8863);
   U9817 : AOI22_X1 port map( A1 => n8752, A2 => n5142, B1 => n8753, B2 => 
                           n5143, ZN => n8861);
   U9818 : AOI22_X1 port map( A1 => n8754, A2 => n5144, B1 => n8755, B2 => 
                           n5145, ZN => n8860);
   U9819 : NAND3_X1 port map( A1 => n8864, A2 => n8865, A3 => n8866, ZN => 
                           n12356);
   U9820 : AOI221_X1 port map( B1 => n8749, B2 => n5149, C1 => n185, C2 => 
                           MEM_IN(28), A => n8867, ZN => n8866);
   U9821 : OAI22_X1 port map( A1 => n10993, A2 => n277, B1 => n5151, B2 => n134
                           , ZN => n8867);
   U9822 : AOI22_X1 port map( A1 => n8752, A2 => n5152, B1 => n8753, B2 => 
                           n5153, ZN => n8865);
   U9823 : AOI22_X1 port map( A1 => n8754, A2 => n5154, B1 => n8755, B2 => 
                           n5155, ZN => n8864);
   U9824 : NAND3_X1 port map( A1 => n8868, A2 => n8869, A3 => n8870, ZN => 
                           n12355);
   U9825 : AOI221_X1 port map( B1 => n8749, B2 => n5159, C1 => n185, C2 => 
                           MEM_IN(29), A => n8871, ZN => n8870);
   U9826 : OAI22_X1 port map( A1 => n10992, A2 => n277, B1 => n5161, B2 => n134
                           , ZN => n8871);
   U9827 : AOI22_X1 port map( A1 => n8752, A2 => n5162, B1 => n8753, B2 => 
                           n5163, ZN => n8869);
   U9828 : AOI22_X1 port map( A1 => n8754, A2 => n5164, B1 => n8755, B2 => 
                           n5165, ZN => n8868);
   U9829 : NAND3_X1 port map( A1 => n8872, A2 => n8873, A3 => n8874, ZN => 
                           n12354);
   U9830 : AOI221_X1 port map( B1 => n8749, B2 => n5169, C1 => n185, C2 => 
                           MEM_IN(30), A => n8875, ZN => n8874);
   U9831 : OAI22_X1 port map( A1 => n10991, A2 => n277, B1 => n5171, B2 => n134
                           , ZN => n8875);
   U9832 : AOI22_X1 port map( A1 => n8752, A2 => n5172, B1 => n8753, B2 => 
                           n5173, ZN => n8873);
   U9833 : AOI22_X1 port map( A1 => n8754, A2 => n5174, B1 => n8755, B2 => 
                           n5175, ZN => n8872);
   U9834 : NAND3_X1 port map( A1 => n8876, A2 => n8877, A3 => n8878, ZN => 
                           n12353);
   U9835 : AOI221_X1 port map( B1 => n8749, B2 => n5179, C1 => n185, C2 => 
                           MEM_IN(31), A => n8879, ZN => n8878);
   U9836 : OAI22_X1 port map( A1 => n10990, A2 => n277, B1 => n5181, B2 => n134
                           , ZN => n8879);
   U9837 : INV_X1 port map( A => n8883, ZN => n8882);
   U9838 : AOI22_X1 port map( A1 => n8752, A2 => n5191, B1 => n8753, B2 => 
                           n5192, ZN => n8877);
   U9839 : AOI22_X1 port map( A1 => n8754, A2 => n5195, B1 => n8755, B2 => 
                           n5196, ZN => n8876);
   U9840 : OAI22_X1 port map( A1 => n8883, A2 => n8881, B1 => n208, B2 => n276,
                           ZN => n8885);
   U9841 : NAND3_X1 port map( A1 => n208, A2 => n277, A3 => n7857, ZN => n8881)
                           ;
   U9842 : INV_X1 port map( A => n8880, ZN => n7857);
   U9843 : OAI22_X1 port map( A1 => n4786, A2 => n8887, B1 => n8888, B2 => 
                           n5204, ZN => n8751);
   U9844 : NOR2_X1 port map( A1 => n8880, A2 => n8883, ZN => n8888);
   U9845 : NAND2_X1 port map( A1 => n8889, A2 => n8447, ZN => n8880);
   U9846 : INV_X1 port map( A => n8890, ZN => n8447);
   U9847 : AOI211_X1 port map( C1 => n8891, C2 => n5207, A => n8892, B => RESET
                           , ZN => n8887);
   U9848 : INV_X1 port map( A => n8884, ZN => n8892);
   U9849 : AOI21_X1 port map( B1 => n8890, B2 => n5206, A => n8886, ZN => n8884
                           );
   U9850 : NAND2_X1 port map( A1 => n8299, A2 => n8303, ZN => n8890);
   U9851 : AND2_X1 port map( A1 => n8155, A2 => n8006, ZN => n8299);
   U9852 : NAND2_X1 port map( A1 => n8893, A2 => n8894, ZN => n8883);
   U9853 : NOR2_X1 port map( A1 => n8006, A2 => n4787, ZN => n8444);
   U9854 : NAND2_X1 port map( A1 => n8895, A2 => n5215, ZN => n8006);
   U9855 : NAND3_X1 port map( A1 => n8896, A2 => n8897, A3 => n8898, ZN => 
                           n12352);
   U9856 : AOI221_X1 port map( B1 => n8899, B2 => n4863, C1 => n178, C2 => 
                           MEM_IN(0), A => n8900, ZN => n8898);
   U9857 : OAI22_X1 port map( A1 => n10989, A2 => n253, B1 => n4867, B2 => n135
                           , ZN => n8900);
   U9858 : AOI22_X1 port map( A1 => n194, A2 => n4869, B1 => n8902, B2 => n4871
                           , ZN => n8897);
   U9859 : AOI22_X1 port map( A1 => n236, A2 => n4873, B1 => n8903, B2 => n4875
                           , ZN => n8896);
   U9860 : NAND3_X1 port map( A1 => n8904, A2 => n8905, A3 => n8906, ZN => 
                           n12351);
   U9861 : AOI221_X1 port map( B1 => n8899, B2 => n4879, C1 => n178, C2 => 
                           MEM_IN(1), A => n8907, ZN => n8906);
   U9862 : OAI22_X1 port map( A1 => n10988, A2 => n253, B1 => n4881, B2 => n135
                           , ZN => n8907);
   U9863 : AOI22_X1 port map( A1 => n194, A2 => n4882, B1 => n8902, B2 => n4883
                           , ZN => n8905);
   U9864 : AOI22_X1 port map( A1 => n236, A2 => n4884, B1 => n8903, B2 => n4885
                           , ZN => n8904);
   U9865 : NAND3_X1 port map( A1 => n8908, A2 => n8909, A3 => n8910, ZN => 
                           n12350);
   U9866 : AOI221_X1 port map( B1 => n8899, B2 => n4889, C1 => n178, C2 => 
                           MEM_IN(2), A => n8911, ZN => n8910);
   U9867 : OAI22_X1 port map( A1 => n10987, A2 => n253, B1 => n4891, B2 => n135
                           , ZN => n8911);
   U9868 : AOI22_X1 port map( A1 => n194, A2 => n4892, B1 => n8902, B2 => n4893
                           , ZN => n8909);
   U9869 : AOI22_X1 port map( A1 => n236, A2 => n4894, B1 => n8903, B2 => n4895
                           , ZN => n8908);
   U9870 : NAND3_X1 port map( A1 => n8912, A2 => n8913, A3 => n8914, ZN => 
                           n12349);
   U9871 : AOI221_X1 port map( B1 => n8899, B2 => n4899, C1 => n178, C2 => 
                           MEM_IN(3), A => n8915, ZN => n8914);
   U9872 : OAI22_X1 port map( A1 => n10986, A2 => n253, B1 => n4901, B2 => n135
                           , ZN => n8915);
   U9873 : AOI22_X1 port map( A1 => n194, A2 => n4902, B1 => n8902, B2 => n4903
                           , ZN => n8913);
   U9874 : AOI22_X1 port map( A1 => n236, A2 => n4904, B1 => n8903, B2 => n4905
                           , ZN => n8912);
   U9875 : NAND3_X1 port map( A1 => n8916, A2 => n8917, A3 => n8918, ZN => 
                           n12348);
   U9876 : AOI221_X1 port map( B1 => n8899, B2 => n4909, C1 => n178, C2 => 
                           MEM_IN(4), A => n8919, ZN => n8918);
   U9877 : OAI22_X1 port map( A1 => n10985, A2 => n253, B1 => n4911, B2 => n135
                           , ZN => n8919);
   U9878 : AOI22_X1 port map( A1 => n194, A2 => n4912, B1 => n8902, B2 => n4913
                           , ZN => n8917);
   U9879 : AOI22_X1 port map( A1 => n236, A2 => n4914, B1 => n8903, B2 => n4915
                           , ZN => n8916);
   U9880 : NAND3_X1 port map( A1 => n8920, A2 => n8921, A3 => n8922, ZN => 
                           n12347);
   U9881 : AOI221_X1 port map( B1 => n8899, B2 => n4919, C1 => n178, C2 => 
                           MEM_IN(5), A => n8923, ZN => n8922);
   U9882 : OAI22_X1 port map( A1 => n10984, A2 => n253, B1 => n4921, B2 => n135
                           , ZN => n8923);
   U9883 : AOI22_X1 port map( A1 => n194, A2 => n4922, B1 => n8902, B2 => n4923
                           , ZN => n8921);
   U9884 : AOI22_X1 port map( A1 => n236, A2 => n4924, B1 => n8903, B2 => n4925
                           , ZN => n8920);
   U9885 : NAND3_X1 port map( A1 => n8924, A2 => n8925, A3 => n8926, ZN => 
                           n12346);
   U9886 : AOI221_X1 port map( B1 => n8899, B2 => n4929, C1 => n178, C2 => 
                           MEM_IN(6), A => n8927, ZN => n8926);
   U9887 : OAI22_X1 port map( A1 => n10983, A2 => n253, B1 => n4931, B2 => n135
                           , ZN => n8927);
   U9888 : AOI22_X1 port map( A1 => n194, A2 => n4932, B1 => n8902, B2 => n4933
                           , ZN => n8925);
   U9889 : AOI22_X1 port map( A1 => n236, A2 => n4934, B1 => n8903, B2 => n4935
                           , ZN => n8924);
   U9890 : NAND3_X1 port map( A1 => n8928, A2 => n8929, A3 => n8930, ZN => 
                           n12345);
   U9891 : AOI221_X1 port map( B1 => n8899, B2 => n4939, C1 => n178, C2 => 
                           MEM_IN(7), A => n8931, ZN => n8930);
   U9892 : OAI22_X1 port map( A1 => n10982, A2 => n253, B1 => n4941, B2 => n135
                           , ZN => n8931);
   U9893 : AOI22_X1 port map( A1 => n194, A2 => n4942, B1 => n8902, B2 => n4943
                           , ZN => n8929);
   U9894 : AOI22_X1 port map( A1 => n236, A2 => n4944, B1 => n8903, B2 => n4945
                           , ZN => n8928);
   U9895 : NAND3_X1 port map( A1 => n8932, A2 => n8933, A3 => n8934, ZN => 
                           n12344);
   U9896 : AOI221_X1 port map( B1 => n8899, B2 => n4949, C1 => n178, C2 => 
                           MEM_IN(8), A => n8935, ZN => n8934);
   U9897 : OAI22_X1 port map( A1 => n10981, A2 => n253, B1 => n4951, B2 => n135
                           , ZN => n8935);
   U9898 : AOI22_X1 port map( A1 => n194, A2 => n4952, B1 => n8902, B2 => n4953
                           , ZN => n8933);
   U9899 : AOI22_X1 port map( A1 => n236, A2 => n4954, B1 => n8903, B2 => n4955
                           , ZN => n8932);
   U9900 : NAND3_X1 port map( A1 => n8936, A2 => n8937, A3 => n8938, ZN => 
                           n12343);
   U9901 : AOI221_X1 port map( B1 => n8899, B2 => n4959, C1 => n178, C2 => 
                           MEM_IN(9), A => n8939, ZN => n8938);
   U9902 : OAI22_X1 port map( A1 => n10980, A2 => n253, B1 => n4961, B2 => n135
                           , ZN => n8939);
   U9903 : AOI22_X1 port map( A1 => n194, A2 => n4962, B1 => n8902, B2 => n4963
                           , ZN => n8937);
   U9904 : AOI22_X1 port map( A1 => n236, A2 => n4964, B1 => n8903, B2 => n4965
                           , ZN => n8936);
   U9905 : NAND3_X1 port map( A1 => n8940, A2 => n8941, A3 => n8942, ZN => 
                           n12342);
   U9906 : AOI221_X1 port map( B1 => n8899, B2 => n4969, C1 => n178, C2 => 
                           MEM_IN(10), A => n8943, ZN => n8942);
   U9907 : OAI22_X1 port map( A1 => n10979, A2 => n253, B1 => n4971, B2 => n135
                           , ZN => n8943);
   U9908 : AOI22_X1 port map( A1 => n194, A2 => n4972, B1 => n8902, B2 => n4973
                           , ZN => n8941);
   U9909 : AOI22_X1 port map( A1 => n236, A2 => n4974, B1 => n8903, B2 => n4975
                           , ZN => n8940);
   U9910 : NAND3_X1 port map( A1 => n8944, A2 => n8945, A3 => n8946, ZN => 
                           n12341);
   U9911 : AOI221_X1 port map( B1 => n8899, B2 => n4979, C1 => n178, C2 => 
                           MEM_IN(11), A => n8947, ZN => n8946);
   U9912 : OAI22_X1 port map( A1 => n10978, A2 => n253, B1 => n4981, B2 => n135
                           , ZN => n8947);
   U9913 : AOI22_X1 port map( A1 => n194, A2 => n4982, B1 => n8902, B2 => n4983
                           , ZN => n8945);
   U9914 : AOI22_X1 port map( A1 => n236, A2 => n4984, B1 => n8903, B2 => n4985
                           , ZN => n8944);
   U9915 : NAND3_X1 port map( A1 => n8948, A2 => n8949, A3 => n8950, ZN => 
                           n12340);
   U9916 : AOI221_X1 port map( B1 => n8899, B2 => n4989, C1 => n178, C2 => 
                           MEM_IN(12), A => n8951, ZN => n8950);
   U9917 : OAI22_X1 port map( A1 => n10977, A2 => n253, B1 => n4991, B2 => n135
                           , ZN => n8951);
   U9918 : AOI22_X1 port map( A1 => n194, A2 => n4992, B1 => n8902, B2 => n4993
                           , ZN => n8949);
   U9919 : AOI22_X1 port map( A1 => n236, A2 => n4994, B1 => n8903, B2 => n4995
                           , ZN => n8948);
   U9920 : NAND3_X1 port map( A1 => n8952, A2 => n8953, A3 => n8954, ZN => 
                           n12339);
   U9921 : AOI221_X1 port map( B1 => n8899, B2 => n4999, C1 => n178, C2 => 
                           MEM_IN(13), A => n8955, ZN => n8954);
   U9922 : OAI22_X1 port map( A1 => n10976, A2 => n253, B1 => n5001, B2 => n135
                           , ZN => n8955);
   U9923 : AOI22_X1 port map( A1 => n194, A2 => n5002, B1 => n8902, B2 => n5003
                           , ZN => n8953);
   U9924 : AOI22_X1 port map( A1 => n236, A2 => n5004, B1 => n8903, B2 => n5005
                           , ZN => n8952);
   U9925 : NAND3_X1 port map( A1 => n8956, A2 => n8957, A3 => n8958, ZN => 
                           n12338);
   U9926 : AOI221_X1 port map( B1 => n8899, B2 => n5009, C1 => n178, C2 => 
                           MEM_IN(14), A => n8959, ZN => n8958);
   U9927 : OAI22_X1 port map( A1 => n10975, A2 => n253, B1 => n5011, B2 => n135
                           , ZN => n8959);
   U9928 : AOI22_X1 port map( A1 => n194, A2 => n5012, B1 => n8902, B2 => n5013
                           , ZN => n8957);
   U9929 : AOI22_X1 port map( A1 => n236, A2 => n5014, B1 => n8903, B2 => n5015
                           , ZN => n8956);
   U9930 : NAND3_X1 port map( A1 => n8960, A2 => n8961, A3 => n8962, ZN => 
                           n12337);
   U9931 : AOI221_X1 port map( B1 => n8899, B2 => n5019, C1 => n178, C2 => 
                           MEM_IN(15), A => n8963, ZN => n8962);
   U9932 : OAI22_X1 port map( A1 => n10974, A2 => n253, B1 => n5021, B2 => n135
                           , ZN => n8963);
   U9933 : AOI22_X1 port map( A1 => n194, A2 => n5022, B1 => n8902, B2 => n5023
                           , ZN => n8961);
   U9934 : AOI22_X1 port map( A1 => n236, A2 => n5024, B1 => n8903, B2 => n5025
                           , ZN => n8960);
   U9935 : NAND3_X1 port map( A1 => n8964, A2 => n8965, A3 => n8966, ZN => 
                           n12336);
   U9936 : AOI221_X1 port map( B1 => n8899, B2 => n5029, C1 => n178, C2 => 
                           MEM_IN(16), A => n8967, ZN => n8966);
   U9937 : OAI22_X1 port map( A1 => n10973, A2 => n253, B1 => n5031, B2 => n135
                           , ZN => n8967);
   U9938 : AOI22_X1 port map( A1 => n194, A2 => n5032, B1 => n8902, B2 => n5033
                           , ZN => n8965);
   U9939 : AOI22_X1 port map( A1 => n236, A2 => n5034, B1 => n8903, B2 => n5035
                           , ZN => n8964);
   U9940 : NAND3_X1 port map( A1 => n8968, A2 => n8969, A3 => n8970, ZN => 
                           n12335);
   U9941 : AOI221_X1 port map( B1 => n8899, B2 => n5039, C1 => n178, C2 => 
                           MEM_IN(17), A => n8971, ZN => n8970);
   U9942 : OAI22_X1 port map( A1 => n10972, A2 => n253, B1 => n5041, B2 => n135
                           , ZN => n8971);
   U9943 : AOI22_X1 port map( A1 => n194, A2 => n5042, B1 => n8902, B2 => n5043
                           , ZN => n8969);
   U9944 : AOI22_X1 port map( A1 => n236, A2 => n5044, B1 => n8903, B2 => n5045
                           , ZN => n8968);
   U9945 : NAND3_X1 port map( A1 => n8972, A2 => n8973, A3 => n8974, ZN => 
                           n12334);
   U9946 : AOI221_X1 port map( B1 => n8899, B2 => n5049, C1 => n178, C2 => 
                           MEM_IN(18), A => n8975, ZN => n8974);
   U9947 : OAI22_X1 port map( A1 => n10971, A2 => n253, B1 => n5051, B2 => n135
                           , ZN => n8975);
   U9948 : AOI22_X1 port map( A1 => n194, A2 => n5052, B1 => n8902, B2 => n5053
                           , ZN => n8973);
   U9949 : AOI22_X1 port map( A1 => n236, A2 => n5054, B1 => n8903, B2 => n5055
                           , ZN => n8972);
   U9950 : NAND3_X1 port map( A1 => n8976, A2 => n8977, A3 => n8978, ZN => 
                           n12333);
   U9951 : AOI221_X1 port map( B1 => n8899, B2 => n5059, C1 => n178, C2 => 
                           MEM_IN(19), A => n8979, ZN => n8978);
   U9952 : OAI22_X1 port map( A1 => n10970, A2 => n253, B1 => n5061, B2 => n135
                           , ZN => n8979);
   U9953 : AOI22_X1 port map( A1 => n194, A2 => n5062, B1 => n8902, B2 => n5063
                           , ZN => n8977);
   U9954 : AOI22_X1 port map( A1 => n236, A2 => n5064, B1 => n8903, B2 => n5065
                           , ZN => n8976);
   U9955 : NAND3_X1 port map( A1 => n8980, A2 => n8981, A3 => n8982, ZN => 
                           n12332);
   U9956 : AOI221_X1 port map( B1 => n8899, B2 => n5069, C1 => n178, C2 => 
                           MEM_IN(20), A => n8983, ZN => n8982);
   U9957 : OAI22_X1 port map( A1 => n10969, A2 => n253, B1 => n5071, B2 => n135
                           , ZN => n8983);
   U9958 : AOI22_X1 port map( A1 => n194, A2 => n5072, B1 => n8902, B2 => n5073
                           , ZN => n8981);
   U9959 : AOI22_X1 port map( A1 => n236, A2 => n5074, B1 => n8903, B2 => n5075
                           , ZN => n8980);
   U9960 : NAND3_X1 port map( A1 => n8984, A2 => n8985, A3 => n8986, ZN => 
                           n12331);
   U9961 : AOI221_X1 port map( B1 => n8899, B2 => n5079, C1 => n178, C2 => 
                           MEM_IN(21), A => n8987, ZN => n8986);
   U9962 : OAI22_X1 port map( A1 => n10968, A2 => n253, B1 => n5081, B2 => n135
                           , ZN => n8987);
   U9963 : AOI22_X1 port map( A1 => n194, A2 => n5082, B1 => n8902, B2 => n5083
                           , ZN => n8985);
   U9964 : AOI22_X1 port map( A1 => n236, A2 => n5084, B1 => n8903, B2 => n5085
                           , ZN => n8984);
   U9965 : NAND3_X1 port map( A1 => n8988, A2 => n8989, A3 => n8990, ZN => 
                           n12330);
   U9966 : AOI221_X1 port map( B1 => n8899, B2 => n5089, C1 => n178, C2 => 
                           MEM_IN(22), A => n8991, ZN => n8990);
   U9967 : OAI22_X1 port map( A1 => n10967, A2 => n253, B1 => n5091, B2 => n135
                           , ZN => n8991);
   U9968 : AOI22_X1 port map( A1 => n194, A2 => n5092, B1 => n8902, B2 => n5093
                           , ZN => n8989);
   U9969 : AOI22_X1 port map( A1 => n236, A2 => n5094, B1 => n8903, B2 => n5095
                           , ZN => n8988);
   U9970 : NAND3_X1 port map( A1 => n8992, A2 => n8993, A3 => n8994, ZN => 
                           n12329);
   U9971 : AOI221_X1 port map( B1 => n8899, B2 => n5099, C1 => n178, C2 => 
                           MEM_IN(23), A => n8995, ZN => n8994);
   U9972 : OAI22_X1 port map( A1 => n10966, A2 => n253, B1 => n5101, B2 => n135
                           , ZN => n8995);
   U9973 : AOI22_X1 port map( A1 => n194, A2 => n5102, B1 => n8902, B2 => n5103
                           , ZN => n8993);
   U9974 : AOI22_X1 port map( A1 => n236, A2 => n5104, B1 => n8903, B2 => n5105
                           , ZN => n8992);
   U9975 : NAND3_X1 port map( A1 => n8996, A2 => n8997, A3 => n8998, ZN => 
                           n12328);
   U9976 : AOI221_X1 port map( B1 => n8899, B2 => n5109, C1 => n178, C2 => 
                           MEM_IN(24), A => n8999, ZN => n8998);
   U9977 : OAI22_X1 port map( A1 => n10965, A2 => n253, B1 => n5111, B2 => n135
                           , ZN => n8999);
   U9978 : AOI22_X1 port map( A1 => n194, A2 => n5112, B1 => n8902, B2 => n5113
                           , ZN => n8997);
   U9979 : AOI22_X1 port map( A1 => n236, A2 => n5114, B1 => n8903, B2 => n5115
                           , ZN => n8996);
   U9980 : NAND3_X1 port map( A1 => n9000, A2 => n9001, A3 => n9002, ZN => 
                           n12327);
   U9981 : AOI221_X1 port map( B1 => n8899, B2 => n5119, C1 => n178, C2 => 
                           MEM_IN(25), A => n9003, ZN => n9002);
   U9982 : OAI22_X1 port map( A1 => n10964, A2 => n253, B1 => n5121, B2 => n135
                           , ZN => n9003);
   U9983 : AOI22_X1 port map( A1 => n194, A2 => n5122, B1 => n8902, B2 => n5123
                           , ZN => n9001);
   U9984 : AOI22_X1 port map( A1 => n236, A2 => n5124, B1 => n8903, B2 => n5125
                           , ZN => n9000);
   U9985 : NAND3_X1 port map( A1 => n9004, A2 => n9005, A3 => n9006, ZN => 
                           n12326);
   U9986 : AOI221_X1 port map( B1 => n8899, B2 => n5129, C1 => n178, C2 => 
                           MEM_IN(26), A => n9007, ZN => n9006);
   U9987 : OAI22_X1 port map( A1 => n10963, A2 => n253, B1 => n5131, B2 => n135
                           , ZN => n9007);
   U9988 : AOI22_X1 port map( A1 => n194, A2 => n5132, B1 => n8902, B2 => n5133
                           , ZN => n9005);
   U9989 : AOI22_X1 port map( A1 => n236, A2 => n5134, B1 => n8903, B2 => n5135
                           , ZN => n9004);
   U9990 : NAND3_X1 port map( A1 => n9008, A2 => n9009, A3 => n9010, ZN => 
                           n12325);
   U9991 : AOI221_X1 port map( B1 => n8899, B2 => n5139, C1 => n178, C2 => 
                           MEM_IN(27), A => n9011, ZN => n9010);
   U9992 : OAI22_X1 port map( A1 => n10962, A2 => n253, B1 => n5141, B2 => n135
                           , ZN => n9011);
   U9993 : AOI22_X1 port map( A1 => n194, A2 => n5142, B1 => n8902, B2 => n5143
                           , ZN => n9009);
   U9994 : AOI22_X1 port map( A1 => n236, A2 => n5144, B1 => n8903, B2 => n5145
                           , ZN => n9008);
   U9995 : NAND3_X1 port map( A1 => n9012, A2 => n9013, A3 => n9014, ZN => 
                           n12324);
   U9996 : AOI221_X1 port map( B1 => n8899, B2 => n5149, C1 => n178, C2 => 
                           MEM_IN(28), A => n9015, ZN => n9014);
   U9997 : OAI22_X1 port map( A1 => n10961, A2 => n253, B1 => n5151, B2 => n135
                           , ZN => n9015);
   U9998 : AOI22_X1 port map( A1 => n194, A2 => n5152, B1 => n8902, B2 => n5153
                           , ZN => n9013);
   U9999 : AOI22_X1 port map( A1 => n236, A2 => n5154, B1 => n8903, B2 => n5155
                           , ZN => n9012);
   U10000 : NAND3_X1 port map( A1 => n9016, A2 => n9017, A3 => n9018, ZN => 
                           n12323);
   U10001 : AOI221_X1 port map( B1 => n8899, B2 => n5159, C1 => n178, C2 => 
                           MEM_IN(29), A => n9019, ZN => n9018);
   U10002 : OAI22_X1 port map( A1 => n10960, A2 => n253, B1 => n5161, B2 => 
                           n135, ZN => n9019);
   U10003 : AOI22_X1 port map( A1 => n194, A2 => n5162, B1 => n8902, B2 => 
                           n5163, ZN => n9017);
   U10004 : AOI22_X1 port map( A1 => n236, A2 => n5164, B1 => n8903, B2 => 
                           n5165, ZN => n9016);
   U10005 : NAND3_X1 port map( A1 => n9020, A2 => n9021, A3 => n9022, ZN => 
                           n12322);
   U10006 : AOI221_X1 port map( B1 => n8899, B2 => n5169, C1 => n178, C2 => 
                           MEM_IN(30), A => n9023, ZN => n9022);
   U10007 : OAI22_X1 port map( A1 => n10959, A2 => n253, B1 => n5171, B2 => 
                           n135, ZN => n9023);
   U10008 : AOI22_X1 port map( A1 => n194, A2 => n5172, B1 => n8902, B2 => 
                           n5173, ZN => n9021);
   U10009 : AOI22_X1 port map( A1 => n236, A2 => n5174, B1 => n8903, B2 => 
                           n5175, ZN => n9020);
   U10010 : NAND3_X1 port map( A1 => n9024, A2 => n9025, A3 => n9026, ZN => 
                           n12321);
   U10011 : AOI221_X1 port map( B1 => n8899, B2 => n5179, C1 => n178, C2 => 
                           MEM_IN(31), A => n9027, ZN => n9026);
   U10012 : OAI22_X1 port map( A1 => n10958, A2 => n253, B1 => n5181, B2 => 
                           n135, ZN => n9027);
   U10013 : AOI22_X1 port map( A1 => n194, A2 => n5191, B1 => n8902, B2 => 
                           n5192, ZN => n9025);
   U10014 : AOI22_X1 port map( A1 => n236, A2 => n5195, B1 => n8903, B2 => 
                           n5196, ZN => n9024);
   U10015 : INV_X1 port map( A => n9034, ZN => n9032);
   U10016 : AOI22_X1 port map( A1 => n9030, A2 => n9037, B1 => n4841, B2 => 
                           n253, ZN => n9034);
   U10017 : INV_X1 port map( A => n9029, ZN => n9037);
   U10018 : NAND3_X1 port map( A1 => n208, A2 => n253, A3 => n8005, ZN => n9029
                           );
   U10019 : INV_X1 port map( A => n9028, ZN => n8005);
   U10020 : OAI22_X1 port map( A1 => n9038, A2 => n4786, B1 => n9039, B2 => 
                           n5204, ZN => n8901);
   U10021 : NOR2_X1 port map( A1 => n9028, A2 => n9040, ZN => n9039);
   U10022 : NAND4_X1 port map( A1 => n8889, A2 => n8894, A3 => n8303, A4 => 
                           n8155, ZN => n9028);
   U10023 : NOR4_X1 port map( A1 => n9041, A2 => n8886, A3 => RESET, A4 => 
                           n9042, ZN => n9038);
   U10024 : OAI211_X1 port map( C1 => n7855, C2 => n9043, A => n8586, B => 
                           n8735, ZN => n9041);
   U10025 : INV_X1 port map( A => n8593, ZN => n8586);
   U10026 : NOR2_X1 port map( A1 => n8155, A2 => n4787, ZN => n8593);
   U10027 : INV_X1 port map( A => n5365, ZN => n7855);
   U10028 : INV_X1 port map( A => n9040, ZN => n9030);
   U10029 : NAND2_X1 port map( A1 => n9044, A2 => n9045, ZN => n9040);
   U10030 : NAND2_X1 port map( A1 => n8895, A2 => n5372, ZN => n8155);
   U10031 : NAND3_X1 port map( A1 => n9046, A2 => n9047, A3 => n9048, ZN => 
                           n12320);
   U10032 : AOI221_X1 port map( B1 => n9049, B2 => n4863, C1 => n179, C2 => 
                           MEM_IN(0), A => n9050, ZN => n9048);
   U10033 : OAI22_X1 port map( A1 => n10957, A2 => n279, B1 => n4867, B2 => 
                           n132, ZN => n9050);
   U10034 : AOI22_X1 port map( A1 => n9052, A2 => n4869, B1 => n9053, B2 => 
                           n4871, ZN => n9047);
   U10035 : AOI22_X1 port map( A1 => n9054, A2 => n4873, B1 => n9055, B2 => 
                           n4875, ZN => n9046);
   U10036 : NAND3_X1 port map( A1 => n9056, A2 => n9057, A3 => n9058, ZN => 
                           n12319);
   U10037 : AOI221_X1 port map( B1 => n9049, B2 => n4879, C1 => n179, C2 => 
                           MEM_IN(1), A => n9059, ZN => n9058);
   U10038 : OAI22_X1 port map( A1 => n10956, A2 => n279, B1 => n4881, B2 => 
                           n132, ZN => n9059);
   U10039 : AOI22_X1 port map( A1 => n9052, A2 => n4882, B1 => n9053, B2 => 
                           n4883, ZN => n9057);
   U10040 : AOI22_X1 port map( A1 => n9054, A2 => n4884, B1 => n9055, B2 => 
                           n4885, ZN => n9056);
   U10041 : NAND3_X1 port map( A1 => n9060, A2 => n9061, A3 => n9062, ZN => 
                           n12318);
   U10042 : AOI221_X1 port map( B1 => n9049, B2 => n4889, C1 => n179, C2 => 
                           MEM_IN(2), A => n9063, ZN => n9062);
   U10043 : OAI22_X1 port map( A1 => n10955, A2 => n279, B1 => n4891, B2 => 
                           n132, ZN => n9063);
   U10044 : AOI22_X1 port map( A1 => n9052, A2 => n4892, B1 => n9053, B2 => 
                           n4893, ZN => n9061);
   U10045 : AOI22_X1 port map( A1 => n9054, A2 => n4894, B1 => n9055, B2 => 
                           n4895, ZN => n9060);
   U10046 : NAND3_X1 port map( A1 => n9064, A2 => n9065, A3 => n9066, ZN => 
                           n12317);
   U10047 : AOI221_X1 port map( B1 => n9049, B2 => n4899, C1 => n179, C2 => 
                           MEM_IN(3), A => n9067, ZN => n9066);
   U10048 : OAI22_X1 port map( A1 => n10954, A2 => n279, B1 => n4901, B2 => 
                           n132, ZN => n9067);
   U10049 : AOI22_X1 port map( A1 => n9052, A2 => n4902, B1 => n9053, B2 => 
                           n4903, ZN => n9065);
   U10050 : AOI22_X1 port map( A1 => n9054, A2 => n4904, B1 => n9055, B2 => 
                           n4905, ZN => n9064);
   U10051 : NAND3_X1 port map( A1 => n9068, A2 => n9069, A3 => n9070, ZN => 
                           n12316);
   U10052 : AOI221_X1 port map( B1 => n9049, B2 => n4909, C1 => n179, C2 => 
                           MEM_IN(4), A => n9071, ZN => n9070);
   U10053 : OAI22_X1 port map( A1 => n10953, A2 => n279, B1 => n4911, B2 => 
                           n132, ZN => n9071);
   U10054 : AOI22_X1 port map( A1 => n9052, A2 => n4912, B1 => n9053, B2 => 
                           n4913, ZN => n9069);
   U10055 : AOI22_X1 port map( A1 => n9054, A2 => n4914, B1 => n9055, B2 => 
                           n4915, ZN => n9068);
   U10056 : NAND3_X1 port map( A1 => n9072, A2 => n9073, A3 => n9074, ZN => 
                           n12315);
   U10057 : AOI221_X1 port map( B1 => n9049, B2 => n4919, C1 => n179, C2 => 
                           MEM_IN(5), A => n9075, ZN => n9074);
   U10058 : OAI22_X1 port map( A1 => n10952, A2 => n279, B1 => n4921, B2 => 
                           n132, ZN => n9075);
   U10059 : AOI22_X1 port map( A1 => n9052, A2 => n4922, B1 => n9053, B2 => 
                           n4923, ZN => n9073);
   U10060 : AOI22_X1 port map( A1 => n9054, A2 => n4924, B1 => n9055, B2 => 
                           n4925, ZN => n9072);
   U10061 : NAND3_X1 port map( A1 => n9076, A2 => n9077, A3 => n9078, ZN => 
                           n12314);
   U10062 : AOI221_X1 port map( B1 => n9049, B2 => n4929, C1 => n179, C2 => 
                           MEM_IN(6), A => n9079, ZN => n9078);
   U10063 : OAI22_X1 port map( A1 => n10951, A2 => n279, B1 => n4931, B2 => 
                           n132, ZN => n9079);
   U10064 : AOI22_X1 port map( A1 => n9052, A2 => n4932, B1 => n9053, B2 => 
                           n4933, ZN => n9077);
   U10065 : AOI22_X1 port map( A1 => n9054, A2 => n4934, B1 => n9055, B2 => 
                           n4935, ZN => n9076);
   U10066 : NAND3_X1 port map( A1 => n9080, A2 => n9081, A3 => n9082, ZN => 
                           n12313);
   U10067 : AOI221_X1 port map( B1 => n9049, B2 => n4939, C1 => n179, C2 => 
                           MEM_IN(7), A => n9083, ZN => n9082);
   U10068 : OAI22_X1 port map( A1 => n10950, A2 => n279, B1 => n4941, B2 => 
                           n132, ZN => n9083);
   U10069 : AOI22_X1 port map( A1 => n9052, A2 => n4942, B1 => n9053, B2 => 
                           n4943, ZN => n9081);
   U10070 : AOI22_X1 port map( A1 => n9054, A2 => n4944, B1 => n9055, B2 => 
                           n4945, ZN => n9080);
   U10071 : NAND3_X1 port map( A1 => n9084, A2 => n9085, A3 => n9086, ZN => 
                           n12312);
   U10072 : AOI221_X1 port map( B1 => n9049, B2 => n4949, C1 => n179, C2 => 
                           MEM_IN(8), A => n9087, ZN => n9086);
   U10073 : OAI22_X1 port map( A1 => n10949, A2 => n279, B1 => n4951, B2 => 
                           n132, ZN => n9087);
   U10074 : AOI22_X1 port map( A1 => n9052, A2 => n4952, B1 => n9053, B2 => 
                           n4953, ZN => n9085);
   U10075 : AOI22_X1 port map( A1 => n9054, A2 => n4954, B1 => n9055, B2 => 
                           n4955, ZN => n9084);
   U10076 : NAND3_X1 port map( A1 => n9088, A2 => n9089, A3 => n9090, ZN => 
                           n12311);
   U10077 : AOI221_X1 port map( B1 => n9049, B2 => n4959, C1 => n179, C2 => 
                           MEM_IN(9), A => n9091, ZN => n9090);
   U10078 : OAI22_X1 port map( A1 => n10948, A2 => n279, B1 => n4961, B2 => 
                           n132, ZN => n9091);
   U10079 : AOI22_X1 port map( A1 => n9052, A2 => n4962, B1 => n9053, B2 => 
                           n4963, ZN => n9089);
   U10080 : AOI22_X1 port map( A1 => n9054, A2 => n4964, B1 => n9055, B2 => 
                           n4965, ZN => n9088);
   U10081 : NAND3_X1 port map( A1 => n9092, A2 => n9093, A3 => n9094, ZN => 
                           n12310);
   U10082 : AOI221_X1 port map( B1 => n9049, B2 => n4969, C1 => n179, C2 => 
                           MEM_IN(10), A => n9095, ZN => n9094);
   U10083 : OAI22_X1 port map( A1 => n10947, A2 => n279, B1 => n4971, B2 => 
                           n132, ZN => n9095);
   U10084 : AOI22_X1 port map( A1 => n9052, A2 => n4972, B1 => n9053, B2 => 
                           n4973, ZN => n9093);
   U10085 : AOI22_X1 port map( A1 => n9054, A2 => n4974, B1 => n9055, B2 => 
                           n4975, ZN => n9092);
   U10086 : NAND3_X1 port map( A1 => n9096, A2 => n9097, A3 => n9098, ZN => 
                           n12309);
   U10087 : AOI221_X1 port map( B1 => n9049, B2 => n4979, C1 => n179, C2 => 
                           MEM_IN(11), A => n9099, ZN => n9098);
   U10088 : OAI22_X1 port map( A1 => n10946, A2 => n279, B1 => n4981, B2 => 
                           n132, ZN => n9099);
   U10089 : AOI22_X1 port map( A1 => n9052, A2 => n4982, B1 => n9053, B2 => 
                           n4983, ZN => n9097);
   U10090 : AOI22_X1 port map( A1 => n9054, A2 => n4984, B1 => n9055, B2 => 
                           n4985, ZN => n9096);
   U10091 : NAND3_X1 port map( A1 => n9100, A2 => n9101, A3 => n9102, ZN => 
                           n12308);
   U10092 : AOI221_X1 port map( B1 => n9049, B2 => n4989, C1 => n179, C2 => 
                           MEM_IN(12), A => n9103, ZN => n9102);
   U10093 : OAI22_X1 port map( A1 => n10945, A2 => n279, B1 => n4991, B2 => 
                           n132, ZN => n9103);
   U10094 : AOI22_X1 port map( A1 => n9052, A2 => n4992, B1 => n9053, B2 => 
                           n4993, ZN => n9101);
   U10095 : AOI22_X1 port map( A1 => n9054, A2 => n4994, B1 => n9055, B2 => 
                           n4995, ZN => n9100);
   U10096 : NAND3_X1 port map( A1 => n9104, A2 => n9105, A3 => n9106, ZN => 
                           n12307);
   U10097 : AOI221_X1 port map( B1 => n9049, B2 => n4999, C1 => n179, C2 => 
                           MEM_IN(13), A => n9107, ZN => n9106);
   U10098 : OAI22_X1 port map( A1 => n10944, A2 => n279, B1 => n5001, B2 => 
                           n132, ZN => n9107);
   U10099 : AOI22_X1 port map( A1 => n9052, A2 => n5002, B1 => n9053, B2 => 
                           n5003, ZN => n9105);
   U10100 : AOI22_X1 port map( A1 => n9054, A2 => n5004, B1 => n9055, B2 => 
                           n5005, ZN => n9104);
   U10101 : NAND3_X1 port map( A1 => n9108, A2 => n9109, A3 => n9110, ZN => 
                           n12306);
   U10102 : AOI221_X1 port map( B1 => n9049, B2 => n5009, C1 => n179, C2 => 
                           MEM_IN(14), A => n9111, ZN => n9110);
   U10103 : OAI22_X1 port map( A1 => n10943, A2 => n279, B1 => n5011, B2 => 
                           n132, ZN => n9111);
   U10104 : AOI22_X1 port map( A1 => n9052, A2 => n5012, B1 => n9053, B2 => 
                           n5013, ZN => n9109);
   U10105 : AOI22_X1 port map( A1 => n9054, A2 => n5014, B1 => n9055, B2 => 
                           n5015, ZN => n9108);
   U10106 : NAND3_X1 port map( A1 => n9112, A2 => n9113, A3 => n9114, ZN => 
                           n12305);
   U10107 : AOI221_X1 port map( B1 => n9049, B2 => n5019, C1 => n179, C2 => 
                           MEM_IN(15), A => n9115, ZN => n9114);
   U10108 : OAI22_X1 port map( A1 => n10942, A2 => n279, B1 => n5021, B2 => 
                           n132, ZN => n9115);
   U10109 : AOI22_X1 port map( A1 => n9052, A2 => n5022, B1 => n9053, B2 => 
                           n5023, ZN => n9113);
   U10110 : AOI22_X1 port map( A1 => n9054, A2 => n5024, B1 => n9055, B2 => 
                           n5025, ZN => n9112);
   U10111 : NAND3_X1 port map( A1 => n9116, A2 => n9117, A3 => n9118, ZN => 
                           n12304);
   U10112 : AOI221_X1 port map( B1 => n9049, B2 => n5029, C1 => n179, C2 => 
                           MEM_IN(16), A => n9119, ZN => n9118);
   U10113 : OAI22_X1 port map( A1 => n10941, A2 => n279, B1 => n5031, B2 => 
                           n132, ZN => n9119);
   U10114 : AOI22_X1 port map( A1 => n9052, A2 => n5032, B1 => n9053, B2 => 
                           n5033, ZN => n9117);
   U10115 : AOI22_X1 port map( A1 => n9054, A2 => n5034, B1 => n9055, B2 => 
                           n5035, ZN => n9116);
   U10116 : NAND3_X1 port map( A1 => n9120, A2 => n9121, A3 => n9122, ZN => 
                           n12303);
   U10117 : AOI221_X1 port map( B1 => n9049, B2 => n5039, C1 => n179, C2 => 
                           MEM_IN(17), A => n9123, ZN => n9122);
   U10118 : OAI22_X1 port map( A1 => n10940, A2 => n279, B1 => n5041, B2 => 
                           n132, ZN => n9123);
   U10119 : AOI22_X1 port map( A1 => n9052, A2 => n5042, B1 => n9053, B2 => 
                           n5043, ZN => n9121);
   U10120 : AOI22_X1 port map( A1 => n9054, A2 => n5044, B1 => n9055, B2 => 
                           n5045, ZN => n9120);
   U10121 : NAND3_X1 port map( A1 => n9124, A2 => n9125, A3 => n9126, ZN => 
                           n12302);
   U10122 : AOI221_X1 port map( B1 => n9049, B2 => n5049, C1 => n179, C2 => 
                           MEM_IN(18), A => n9127, ZN => n9126);
   U10123 : OAI22_X1 port map( A1 => n10939, A2 => n279, B1 => n5051, B2 => 
                           n132, ZN => n9127);
   U10124 : AOI22_X1 port map( A1 => n9052, A2 => n5052, B1 => n9053, B2 => 
                           n5053, ZN => n9125);
   U10125 : AOI22_X1 port map( A1 => n9054, A2 => n5054, B1 => n9055, B2 => 
                           n5055, ZN => n9124);
   U10126 : NAND3_X1 port map( A1 => n9128, A2 => n9129, A3 => n9130, ZN => 
                           n12301);
   U10127 : AOI221_X1 port map( B1 => n9049, B2 => n5059, C1 => n179, C2 => 
                           MEM_IN(19), A => n9131, ZN => n9130);
   U10128 : OAI22_X1 port map( A1 => n10938, A2 => n279, B1 => n5061, B2 => 
                           n132, ZN => n9131);
   U10129 : AOI22_X1 port map( A1 => n9052, A2 => n5062, B1 => n9053, B2 => 
                           n5063, ZN => n9129);
   U10130 : AOI22_X1 port map( A1 => n9054, A2 => n5064, B1 => n9055, B2 => 
                           n5065, ZN => n9128);
   U10131 : NAND3_X1 port map( A1 => n9132, A2 => n9133, A3 => n9134, ZN => 
                           n12300_port);
   U10132 : AOI221_X1 port map( B1 => n9049, B2 => n5069, C1 => n179, C2 => 
                           MEM_IN(20), A => n9135, ZN => n9134);
   U10133 : OAI22_X1 port map( A1 => n10937, A2 => n279, B1 => n5071, B2 => 
                           n132, ZN => n9135);
   U10134 : AOI22_X1 port map( A1 => n9052, A2 => n5072, B1 => n9053, B2 => 
                           n5073, ZN => n9133);
   U10135 : AOI22_X1 port map( A1 => n9054, A2 => n5074, B1 => n9055, B2 => 
                           n5075, ZN => n9132);
   U10136 : NAND3_X1 port map( A1 => n9136, A2 => n9137, A3 => n9138, ZN => 
                           n12299_port);
   U10137 : AOI221_X1 port map( B1 => n9049, B2 => n5079, C1 => n179, C2 => 
                           MEM_IN(21), A => n9139, ZN => n9138);
   U10138 : OAI22_X1 port map( A1 => n10936, A2 => n279, B1 => n5081, B2 => 
                           n132, ZN => n9139);
   U10139 : AOI22_X1 port map( A1 => n9052, A2 => n5082, B1 => n9053, B2 => 
                           n5083, ZN => n9137);
   U10140 : AOI22_X1 port map( A1 => n9054, A2 => n5084, B1 => n9055, B2 => 
                           n5085, ZN => n9136);
   U10141 : NAND3_X1 port map( A1 => n9140, A2 => n9141, A3 => n9142, ZN => 
                           n12298_port);
   U10142 : AOI221_X1 port map( B1 => n9049, B2 => n5089, C1 => n179, C2 => 
                           MEM_IN(22), A => n9143, ZN => n9142);
   U10143 : OAI22_X1 port map( A1 => n10935, A2 => n279, B1 => n5091, B2 => 
                           n132, ZN => n9143);
   U10144 : AOI22_X1 port map( A1 => n9052, A2 => n5092, B1 => n9053, B2 => 
                           n5093, ZN => n9141);
   U10145 : AOI22_X1 port map( A1 => n9054, A2 => n5094, B1 => n9055, B2 => 
                           n5095, ZN => n9140);
   U10146 : NAND3_X1 port map( A1 => n9144, A2 => n9145, A3 => n9146, ZN => 
                           n12297_port);
   U10147 : AOI221_X1 port map( B1 => n9049, B2 => n5099, C1 => n179, C2 => 
                           MEM_IN(23), A => n9147, ZN => n9146);
   U10148 : OAI22_X1 port map( A1 => n10934, A2 => n279, B1 => n5101, B2 => 
                           n132, ZN => n9147);
   U10149 : AOI22_X1 port map( A1 => n9052, A2 => n5102, B1 => n9053, B2 => 
                           n5103, ZN => n9145);
   U10150 : AOI22_X1 port map( A1 => n9054, A2 => n5104, B1 => n9055, B2 => 
                           n5105, ZN => n9144);
   U10151 : NAND3_X1 port map( A1 => n9148, A2 => n9149, A3 => n9150, ZN => 
                           n12296_port);
   U10152 : AOI221_X1 port map( B1 => n9049, B2 => n5109, C1 => n179, C2 => 
                           MEM_IN(24), A => n9151, ZN => n9150);
   U10153 : OAI22_X1 port map( A1 => n10933, A2 => n279, B1 => n5111, B2 => 
                           n132, ZN => n9151);
   U10154 : AOI22_X1 port map( A1 => n9052, A2 => n5112, B1 => n9053, B2 => 
                           n5113, ZN => n9149);
   U10155 : AOI22_X1 port map( A1 => n9054, A2 => n5114, B1 => n9055, B2 => 
                           n5115, ZN => n9148);
   U10156 : NAND3_X1 port map( A1 => n9152, A2 => n9153, A3 => n9154, ZN => 
                           n12295_port);
   U10157 : AOI221_X1 port map( B1 => n9049, B2 => n5119, C1 => n179, C2 => 
                           MEM_IN(25), A => n9155, ZN => n9154);
   U10158 : OAI22_X1 port map( A1 => n10932, A2 => n279, B1 => n5121, B2 => 
                           n132, ZN => n9155);
   U10159 : AOI22_X1 port map( A1 => n9052, A2 => n5122, B1 => n9053, B2 => 
                           n5123, ZN => n9153);
   U10160 : AOI22_X1 port map( A1 => n9054, A2 => n5124, B1 => n9055, B2 => 
                           n5125, ZN => n9152);
   U10161 : NAND3_X1 port map( A1 => n9156, A2 => n9157, A3 => n9158, ZN => 
                           n12294_port);
   U10162 : AOI221_X1 port map( B1 => n9049, B2 => n5129, C1 => n179, C2 => 
                           MEM_IN(26), A => n9159, ZN => n9158);
   U10163 : OAI22_X1 port map( A1 => n10931, A2 => n279, B1 => n5131, B2 => 
                           n132, ZN => n9159);
   U10164 : AOI22_X1 port map( A1 => n9052, A2 => n5132, B1 => n9053, B2 => 
                           n5133, ZN => n9157);
   U10165 : AOI22_X1 port map( A1 => n9054, A2 => n5134, B1 => n9055, B2 => 
                           n5135, ZN => n9156);
   U10166 : NAND3_X1 port map( A1 => n9160, A2 => n9161, A3 => n9162, ZN => 
                           n12293_port);
   U10167 : AOI221_X1 port map( B1 => n9049, B2 => n5139, C1 => n179, C2 => 
                           MEM_IN(27), A => n9163, ZN => n9162);
   U10168 : OAI22_X1 port map( A1 => n10930, A2 => n279, B1 => n5141, B2 => 
                           n132, ZN => n9163);
   U10169 : AOI22_X1 port map( A1 => n9052, A2 => n5142, B1 => n9053, B2 => 
                           n5143, ZN => n9161);
   U10170 : AOI22_X1 port map( A1 => n9054, A2 => n5144, B1 => n9055, B2 => 
                           n5145, ZN => n9160);
   U10171 : NAND3_X1 port map( A1 => n9164, A2 => n9165, A3 => n9166, ZN => 
                           n12292_port);
   U10172 : AOI221_X1 port map( B1 => n9049, B2 => n5149, C1 => n179, C2 => 
                           MEM_IN(28), A => n9167, ZN => n9166);
   U10173 : OAI22_X1 port map( A1 => n10929, A2 => n279, B1 => n5151, B2 => 
                           n132, ZN => n9167);
   U10174 : AOI22_X1 port map( A1 => n9052, A2 => n5152, B1 => n9053, B2 => 
                           n5153, ZN => n9165);
   U10175 : AOI22_X1 port map( A1 => n9054, A2 => n5154, B1 => n9055, B2 => 
                           n5155, ZN => n9164);
   U10176 : NAND3_X1 port map( A1 => n9168, A2 => n9169, A3 => n9170, ZN => 
                           n12291_port);
   U10177 : AOI221_X1 port map( B1 => n9049, B2 => n5159, C1 => n179, C2 => 
                           MEM_IN(29), A => n9171, ZN => n9170);
   U10178 : OAI22_X1 port map( A1 => n10928, A2 => n279, B1 => n5161, B2 => 
                           n132, ZN => n9171);
   U10179 : AOI22_X1 port map( A1 => n9052, A2 => n5162, B1 => n9053, B2 => 
                           n5163, ZN => n9169);
   U10180 : AOI22_X1 port map( A1 => n9054, A2 => n5164, B1 => n9055, B2 => 
                           n5165, ZN => n9168);
   U10181 : NAND3_X1 port map( A1 => n9172, A2 => n9173, A3 => n9174, ZN => 
                           n12290_port);
   U10182 : AOI221_X1 port map( B1 => n9049, B2 => n5169, C1 => n179, C2 => 
                           MEM_IN(30), A => n9175, ZN => n9174);
   U10183 : OAI22_X1 port map( A1 => n10927, A2 => n279, B1 => n5171, B2 => 
                           n132, ZN => n9175);
   U10184 : AOI22_X1 port map( A1 => n9052, A2 => n5172, B1 => n9053, B2 => 
                           n5173, ZN => n9173);
   U10185 : AOI22_X1 port map( A1 => n9054, A2 => n5174, B1 => n9055, B2 => 
                           n5175, ZN => n9172);
   U10186 : NAND3_X1 port map( A1 => n9176, A2 => n9177, A3 => n9178, ZN => 
                           n12289_port);
   U10187 : AOI221_X1 port map( B1 => n9049, B2 => n5179, C1 => n179, C2 => 
                           MEM_IN(31), A => n9179, ZN => n9178);
   U10188 : OAI22_X1 port map( A1 => n10926, A2 => n279, B1 => n5181, B2 => 
                           n132, ZN => n9179);
   U10189 : INV_X1 port map( A => n9183, ZN => n9182);
   U10190 : INV_X1 port map( A => n8737, ZN => n8735);
   U10191 : AOI22_X1 port map( A1 => n9052, A2 => n5191, B1 => n9053, B2 => 
                           n5192, ZN => n9177);
   U10192 : AOI22_X1 port map( A1 => n9054, A2 => n5195, B1 => n9055, B2 => 
                           n5196, ZN => n9176);
   U10193 : OAI22_X1 port map( A1 => n9183, A2 => n9181, B1 => n208, B2 => n278
                           , ZN => n9184);
   U10194 : NAND3_X1 port map( A1 => n208, A2 => n279, A3 => n8154, ZN => n9181
                           );
   U10195 : INV_X1 port map( A => n9180, ZN => n8154);
   U10196 : OAI22_X1 port map( A1 => n4786, A2 => n9187, B1 => n9188, B2 => 
                           n5204, ZN => n9051);
   U10197 : NOR2_X1 port map( A1 => n9180, A2 => n9183, ZN => n9188);
   U10198 : NAND3_X1 port map( A1 => n8889, A2 => n8303, A3 => n9189, ZN => 
                           n9180);
   U10199 : AOI211_X1 port map( C1 => n8891, C2 => n5522, A => n9190, B => 
                           n8737, ZN => n9187);
   U10200 : NOR2_X1 port map( A1 => n8303, A2 => n4787, ZN => n8737);
   U10201 : NAND2_X1 port map( A1 => n9191, A2 => n9192, ZN => n9183);
   U10202 : NOR2_X1 port map( A1 => n9036, A2 => n8303, ZN => n9035);
   U10203 : NAND2_X1 port map( A1 => n8895, A2 => n5526, ZN => n8303);
   U10204 : NAND3_X1 port map( A1 => n9193, A2 => n9194, A3 => n9195, ZN => 
                           n12288_port);
   U10205 : AOI221_X1 port map( B1 => n9196, B2 => n4863, C1 => n180, C2 => 
                           MEM_IN(0), A => n9197, ZN => n9195);
   U10206 : OAI22_X1 port map( A1 => n10925, A2 => n281, B1 => n4867, B2 => 
                           n133, ZN => n9197);
   U10207 : AOI22_X1 port map( A1 => n9199, A2 => n4869, B1 => n9200, B2 => 
                           n4871, ZN => n9194);
   U10208 : AOI22_X1 port map( A1 => n9201, A2 => n4873, B1 => n9202, B2 => 
                           n4875, ZN => n9193);
   U10209 : NAND3_X1 port map( A1 => n9203, A2 => n9204, A3 => n9205, ZN => 
                           n12287_port);
   U10210 : AOI221_X1 port map( B1 => n9196, B2 => n4879, C1 => n180, C2 => 
                           MEM_IN(1), A => n9206, ZN => n9205);
   U10211 : OAI22_X1 port map( A1 => n10924, A2 => n281, B1 => n4881, B2 => 
                           n133, ZN => n9206);
   U10212 : AOI22_X1 port map( A1 => n9199, A2 => n4882, B1 => n9200, B2 => 
                           n4883, ZN => n9204);
   U10213 : AOI22_X1 port map( A1 => n9201, A2 => n4884, B1 => n9202, B2 => 
                           n4885, ZN => n9203);
   U10214 : NAND3_X1 port map( A1 => n9207, A2 => n9208, A3 => n9209, ZN => 
                           n12286_port);
   U10215 : AOI221_X1 port map( B1 => n9196, B2 => n4889, C1 => n180, C2 => 
                           MEM_IN(2), A => n9210, ZN => n9209);
   U10216 : OAI22_X1 port map( A1 => n10923, A2 => n281, B1 => n4891, B2 => 
                           n133, ZN => n9210);
   U10217 : AOI22_X1 port map( A1 => n9199, A2 => n4892, B1 => n9200, B2 => 
                           n4893, ZN => n9208);
   U10218 : AOI22_X1 port map( A1 => n9201, A2 => n4894, B1 => n9202, B2 => 
                           n4895, ZN => n9207);
   U10219 : NAND3_X1 port map( A1 => n9211, A2 => n9212, A3 => n9213, ZN => 
                           n12285_port);
   U10220 : AOI221_X1 port map( B1 => n9196, B2 => n4899, C1 => n180, C2 => 
                           MEM_IN(3), A => n9214, ZN => n9213);
   U10221 : OAI22_X1 port map( A1 => n10922, A2 => n281, B1 => n4901, B2 => 
                           n133, ZN => n9214);
   U10222 : AOI22_X1 port map( A1 => n9199, A2 => n4902, B1 => n9200, B2 => 
                           n4903, ZN => n9212);
   U10223 : AOI22_X1 port map( A1 => n9201, A2 => n4904, B1 => n9202, B2 => 
                           n4905, ZN => n9211);
   U10224 : NAND3_X1 port map( A1 => n9215, A2 => n9216, A3 => n9217, ZN => 
                           n12284_port);
   U10225 : AOI221_X1 port map( B1 => n9196, B2 => n4909, C1 => n180, C2 => 
                           MEM_IN(4), A => n9218, ZN => n9217);
   U10226 : OAI22_X1 port map( A1 => n10921, A2 => n281, B1 => n4911, B2 => 
                           n133, ZN => n9218);
   U10227 : AOI22_X1 port map( A1 => n9199, A2 => n4912, B1 => n9200, B2 => 
                           n4913, ZN => n9216);
   U10228 : AOI22_X1 port map( A1 => n9201, A2 => n4914, B1 => n9202, B2 => 
                           n4915, ZN => n9215);
   U10229 : NAND3_X1 port map( A1 => n9219, A2 => n9220, A3 => n9221, ZN => 
                           n12283_port);
   U10230 : AOI221_X1 port map( B1 => n9196, B2 => n4919, C1 => n180, C2 => 
                           MEM_IN(5), A => n9222, ZN => n9221);
   U10231 : OAI22_X1 port map( A1 => n10920, A2 => n281, B1 => n4921, B2 => 
                           n133, ZN => n9222);
   U10232 : AOI22_X1 port map( A1 => n9199, A2 => n4922, B1 => n9200, B2 => 
                           n4923, ZN => n9220);
   U10233 : AOI22_X1 port map( A1 => n9201, A2 => n4924, B1 => n9202, B2 => 
                           n4925, ZN => n9219);
   U10234 : NAND3_X1 port map( A1 => n9223, A2 => n9224, A3 => n9225, ZN => 
                           n12282_port);
   U10235 : AOI221_X1 port map( B1 => n9196, B2 => n4929, C1 => n180, C2 => 
                           MEM_IN(6), A => n9226, ZN => n9225);
   U10236 : OAI22_X1 port map( A1 => n10919, A2 => n281, B1 => n4931, B2 => 
                           n133, ZN => n9226);
   U10237 : AOI22_X1 port map( A1 => n9199, A2 => n4932, B1 => n9200, B2 => 
                           n4933, ZN => n9224);
   U10238 : AOI22_X1 port map( A1 => n9201, A2 => n4934, B1 => n9202, B2 => 
                           n4935, ZN => n9223);
   U10239 : NAND3_X1 port map( A1 => n9227, A2 => n9228, A3 => n9229, ZN => 
                           n12281_port);
   U10240 : AOI221_X1 port map( B1 => n9196, B2 => n4939, C1 => n180, C2 => 
                           MEM_IN(7), A => n9230, ZN => n9229);
   U10241 : OAI22_X1 port map( A1 => n10918, A2 => n281, B1 => n4941, B2 => 
                           n133, ZN => n9230);
   U10242 : AOI22_X1 port map( A1 => n9199, A2 => n4942, B1 => n9200, B2 => 
                           n4943, ZN => n9228);
   U10243 : AOI22_X1 port map( A1 => n9201, A2 => n4944, B1 => n9202, B2 => 
                           n4945, ZN => n9227);
   U10244 : NAND3_X1 port map( A1 => n9231, A2 => n9232, A3 => n9233, ZN => 
                           n12280_port);
   U10245 : AOI221_X1 port map( B1 => n9196, B2 => n4949, C1 => n180, C2 => 
                           MEM_IN(8), A => n9234, ZN => n9233);
   U10246 : OAI22_X1 port map( A1 => n10917, A2 => n281, B1 => n4951, B2 => 
                           n133, ZN => n9234);
   U10247 : AOI22_X1 port map( A1 => n9199, A2 => n4952, B1 => n9200, B2 => 
                           n4953, ZN => n9232);
   U10248 : AOI22_X1 port map( A1 => n9201, A2 => n4954, B1 => n9202, B2 => 
                           n4955, ZN => n9231);
   U10249 : NAND3_X1 port map( A1 => n9235, A2 => n9236, A3 => n9237, ZN => 
                           n12279_port);
   U10250 : AOI221_X1 port map( B1 => n9196, B2 => n4959, C1 => n180, C2 => 
                           MEM_IN(9), A => n9238, ZN => n9237);
   U10251 : OAI22_X1 port map( A1 => n10916, A2 => n281, B1 => n4961, B2 => 
                           n133, ZN => n9238);
   U10252 : AOI22_X1 port map( A1 => n9199, A2 => n4962, B1 => n9200, B2 => 
                           n4963, ZN => n9236);
   U10253 : AOI22_X1 port map( A1 => n9201, A2 => n4964, B1 => n9202, B2 => 
                           n4965, ZN => n9235);
   U10254 : NAND3_X1 port map( A1 => n9239, A2 => n9240, A3 => n9241, ZN => 
                           n12278_port);
   U10255 : AOI221_X1 port map( B1 => n9196, B2 => n4969, C1 => n180, C2 => 
                           MEM_IN(10), A => n9242, ZN => n9241);
   U10256 : OAI22_X1 port map( A1 => n10915, A2 => n281, B1 => n4971, B2 => 
                           n133, ZN => n9242);
   U10257 : AOI22_X1 port map( A1 => n9199, A2 => n4972, B1 => n9200, B2 => 
                           n4973, ZN => n9240);
   U10258 : AOI22_X1 port map( A1 => n9201, A2 => n4974, B1 => n9202, B2 => 
                           n4975, ZN => n9239);
   U10259 : NAND3_X1 port map( A1 => n9243, A2 => n9244, A3 => n9245, ZN => 
                           n12277_port);
   U10260 : AOI221_X1 port map( B1 => n9196, B2 => n4979, C1 => n180, C2 => 
                           MEM_IN(11), A => n9246, ZN => n9245);
   U10261 : OAI22_X1 port map( A1 => n10914, A2 => n281, B1 => n4981, B2 => 
                           n133, ZN => n9246);
   U10262 : AOI22_X1 port map( A1 => n9199, A2 => n4982, B1 => n9200, B2 => 
                           n4983, ZN => n9244);
   U10263 : AOI22_X1 port map( A1 => n9201, A2 => n4984, B1 => n9202, B2 => 
                           n4985, ZN => n9243);
   U10264 : NAND3_X1 port map( A1 => n9247, A2 => n9248, A3 => n9249, ZN => 
                           n12276_port);
   U10265 : AOI221_X1 port map( B1 => n9196, B2 => n4989, C1 => n180, C2 => 
                           MEM_IN(12), A => n9250, ZN => n9249);
   U10266 : OAI22_X1 port map( A1 => n10913, A2 => n281, B1 => n4991, B2 => 
                           n133, ZN => n9250);
   U10267 : AOI22_X1 port map( A1 => n9199, A2 => n4992, B1 => n9200, B2 => 
                           n4993, ZN => n9248);
   U10268 : AOI22_X1 port map( A1 => n9201, A2 => n4994, B1 => n9202, B2 => 
                           n4995, ZN => n9247);
   U10269 : NAND3_X1 port map( A1 => n9251, A2 => n9252, A3 => n9253, ZN => 
                           n12275_port);
   U10270 : AOI221_X1 port map( B1 => n9196, B2 => n4999, C1 => n180, C2 => 
                           MEM_IN(13), A => n9254, ZN => n9253);
   U10271 : OAI22_X1 port map( A1 => n10912, A2 => n281, B1 => n5001, B2 => 
                           n133, ZN => n9254);
   U10272 : AOI22_X1 port map( A1 => n9199, A2 => n5002, B1 => n9200, B2 => 
                           n5003, ZN => n9252);
   U10273 : AOI22_X1 port map( A1 => n9201, A2 => n5004, B1 => n9202, B2 => 
                           n5005, ZN => n9251);
   U10274 : NAND3_X1 port map( A1 => n9255, A2 => n9256, A3 => n9257, ZN => 
                           n12274_port);
   U10275 : AOI221_X1 port map( B1 => n9196, B2 => n5009, C1 => n180, C2 => 
                           MEM_IN(14), A => n9258, ZN => n9257);
   U10276 : OAI22_X1 port map( A1 => n10911, A2 => n281, B1 => n5011, B2 => 
                           n133, ZN => n9258);
   U10277 : AOI22_X1 port map( A1 => n9199, A2 => n5012, B1 => n9200, B2 => 
                           n5013, ZN => n9256);
   U10278 : AOI22_X1 port map( A1 => n9201, A2 => n5014, B1 => n9202, B2 => 
                           n5015, ZN => n9255);
   U10279 : NAND3_X1 port map( A1 => n9259, A2 => n9260, A3 => n9261, ZN => 
                           n12273_port);
   U10280 : AOI221_X1 port map( B1 => n9196, B2 => n5019, C1 => n180, C2 => 
                           MEM_IN(15), A => n9262, ZN => n9261);
   U10281 : OAI22_X1 port map( A1 => n10910, A2 => n281, B1 => n5021, B2 => 
                           n133, ZN => n9262);
   U10282 : AOI22_X1 port map( A1 => n9199, A2 => n5022, B1 => n9200, B2 => 
                           n5023, ZN => n9260);
   U10283 : AOI22_X1 port map( A1 => n9201, A2 => n5024, B1 => n9202, B2 => 
                           n5025, ZN => n9259);
   U10284 : NAND3_X1 port map( A1 => n9263, A2 => n9264, A3 => n9265, ZN => 
                           n12272_port);
   U10285 : AOI221_X1 port map( B1 => n9196, B2 => n5029, C1 => n180, C2 => 
                           MEM_IN(16), A => n9266, ZN => n9265);
   U10286 : OAI22_X1 port map( A1 => n10909, A2 => n281, B1 => n5031, B2 => 
                           n133, ZN => n9266);
   U10287 : AOI22_X1 port map( A1 => n9199, A2 => n5032, B1 => n9200, B2 => 
                           n5033, ZN => n9264);
   U10288 : AOI22_X1 port map( A1 => n9201, A2 => n5034, B1 => n9202, B2 => 
                           n5035, ZN => n9263);
   U10289 : NAND3_X1 port map( A1 => n9267, A2 => n9268, A3 => n9269, ZN => 
                           n12271_port);
   U10290 : AOI221_X1 port map( B1 => n9196, B2 => n5039, C1 => n180, C2 => 
                           MEM_IN(17), A => n9270, ZN => n9269);
   U10291 : OAI22_X1 port map( A1 => n10908, A2 => n281, B1 => n5041, B2 => 
                           n133, ZN => n9270);
   U10292 : AOI22_X1 port map( A1 => n9199, A2 => n5042, B1 => n9200, B2 => 
                           n5043, ZN => n9268);
   U10293 : AOI22_X1 port map( A1 => n9201, A2 => n5044, B1 => n9202, B2 => 
                           n5045, ZN => n9267);
   U10294 : NAND3_X1 port map( A1 => n9271, A2 => n9272, A3 => n9273, ZN => 
                           n12270_port);
   U10295 : AOI221_X1 port map( B1 => n9196, B2 => n5049, C1 => n180, C2 => 
                           MEM_IN(18), A => n9274, ZN => n9273);
   U10296 : OAI22_X1 port map( A1 => n10907, A2 => n281, B1 => n5051, B2 => 
                           n133, ZN => n9274);
   U10297 : AOI22_X1 port map( A1 => n9199, A2 => n5052, B1 => n9200, B2 => 
                           n5053, ZN => n9272);
   U10298 : AOI22_X1 port map( A1 => n9201, A2 => n5054, B1 => n9202, B2 => 
                           n5055, ZN => n9271);
   U10299 : NAND3_X1 port map( A1 => n9275, A2 => n9276, A3 => n9277, ZN => 
                           n12269_port);
   U10300 : AOI221_X1 port map( B1 => n9196, B2 => n5059, C1 => n180, C2 => 
                           MEM_IN(19), A => n9278, ZN => n9277);
   U10301 : OAI22_X1 port map( A1 => n10906, A2 => n281, B1 => n5061, B2 => 
                           n133, ZN => n9278);
   U10302 : AOI22_X1 port map( A1 => n9199, A2 => n5062, B1 => n9200, B2 => 
                           n5063, ZN => n9276);
   U10303 : AOI22_X1 port map( A1 => n9201, A2 => n5064, B1 => n9202, B2 => 
                           n5065, ZN => n9275);
   U10304 : NAND3_X1 port map( A1 => n9279, A2 => n9280, A3 => n9281, ZN => 
                           n12268_port);
   U10305 : AOI221_X1 port map( B1 => n9196, B2 => n5069, C1 => n180, C2 => 
                           MEM_IN(20), A => n9282, ZN => n9281);
   U10306 : OAI22_X1 port map( A1 => n10905, A2 => n281, B1 => n5071, B2 => 
                           n133, ZN => n9282);
   U10307 : AOI22_X1 port map( A1 => n9199, A2 => n5072, B1 => n9200, B2 => 
                           n5073, ZN => n9280);
   U10308 : AOI22_X1 port map( A1 => n9201, A2 => n5074, B1 => n9202, B2 => 
                           n5075, ZN => n9279);
   U10309 : NAND3_X1 port map( A1 => n9283, A2 => n9284, A3 => n9285, ZN => 
                           n12267_port);
   U10310 : AOI221_X1 port map( B1 => n9196, B2 => n5079, C1 => n180, C2 => 
                           MEM_IN(21), A => n9286, ZN => n9285);
   U10311 : OAI22_X1 port map( A1 => n10904, A2 => n281, B1 => n5081, B2 => 
                           n133, ZN => n9286);
   U10312 : AOI22_X1 port map( A1 => n9199, A2 => n5082, B1 => n9200, B2 => 
                           n5083, ZN => n9284);
   U10313 : AOI22_X1 port map( A1 => n9201, A2 => n5084, B1 => n9202, B2 => 
                           n5085, ZN => n9283);
   U10314 : NAND3_X1 port map( A1 => n9287, A2 => n9288, A3 => n9289, ZN => 
                           n12266_port);
   U10315 : AOI221_X1 port map( B1 => n9196, B2 => n5089, C1 => n180, C2 => 
                           MEM_IN(22), A => n9290, ZN => n9289);
   U10316 : OAI22_X1 port map( A1 => n10903, A2 => n281, B1 => n5091, B2 => 
                           n133, ZN => n9290);
   U10317 : AOI22_X1 port map( A1 => n9199, A2 => n5092, B1 => n9200, B2 => 
                           n5093, ZN => n9288);
   U10318 : AOI22_X1 port map( A1 => n9201, A2 => n5094, B1 => n9202, B2 => 
                           n5095, ZN => n9287);
   U10319 : NAND3_X1 port map( A1 => n9291, A2 => n9292, A3 => n9293, ZN => 
                           n12265_port);
   U10320 : AOI221_X1 port map( B1 => n9196, B2 => n5099, C1 => n180, C2 => 
                           MEM_IN(23), A => n9294, ZN => n9293);
   U10321 : OAI22_X1 port map( A1 => n10902, A2 => n281, B1 => n5101, B2 => 
                           n133, ZN => n9294);
   U10322 : AOI22_X1 port map( A1 => n9199, A2 => n5102, B1 => n9200, B2 => 
                           n5103, ZN => n9292);
   U10323 : AOI22_X1 port map( A1 => n9201, A2 => n5104, B1 => n9202, B2 => 
                           n5105, ZN => n9291);
   U10324 : NAND3_X1 port map( A1 => n9295, A2 => n9296, A3 => n9297, ZN => 
                           n12264_port);
   U10325 : AOI221_X1 port map( B1 => n9196, B2 => n5109, C1 => n180, C2 => 
                           MEM_IN(24), A => n9298, ZN => n9297);
   U10326 : OAI22_X1 port map( A1 => n10901, A2 => n281, B1 => n5111, B2 => 
                           n133, ZN => n9298);
   U10327 : AOI22_X1 port map( A1 => n9199, A2 => n5112, B1 => n9200, B2 => 
                           n5113, ZN => n9296);
   U10328 : AOI22_X1 port map( A1 => n9201, A2 => n5114, B1 => n9202, B2 => 
                           n5115, ZN => n9295);
   U10329 : NAND3_X1 port map( A1 => n9299, A2 => n9300, A3 => n9301, ZN => 
                           n12263_port);
   U10330 : AOI221_X1 port map( B1 => n9196, B2 => n5119, C1 => n180, C2 => 
                           MEM_IN(25), A => n9302, ZN => n9301);
   U10331 : OAI22_X1 port map( A1 => n10900, A2 => n281, B1 => n5121, B2 => 
                           n133, ZN => n9302);
   U10332 : AOI22_X1 port map( A1 => n9199, A2 => n5122, B1 => n9200, B2 => 
                           n5123, ZN => n9300);
   U10333 : AOI22_X1 port map( A1 => n9201, A2 => n5124, B1 => n9202, B2 => 
                           n5125, ZN => n9299);
   U10334 : NAND3_X1 port map( A1 => n9303, A2 => n9304, A3 => n9305, ZN => 
                           n12262_port);
   U10335 : AOI221_X1 port map( B1 => n9196, B2 => n5129, C1 => n180, C2 => 
                           MEM_IN(26), A => n9306, ZN => n9305);
   U10336 : OAI22_X1 port map( A1 => n10899, A2 => n281, B1 => n5131, B2 => 
                           n133, ZN => n9306);
   U10337 : AOI22_X1 port map( A1 => n9199, A2 => n5132, B1 => n9200, B2 => 
                           n5133, ZN => n9304);
   U10338 : AOI22_X1 port map( A1 => n9201, A2 => n5134, B1 => n9202, B2 => 
                           n5135, ZN => n9303);
   U10339 : NAND3_X1 port map( A1 => n9307, A2 => n9308, A3 => n9309, ZN => 
                           n12261_port);
   U10340 : AOI221_X1 port map( B1 => n9196, B2 => n5139, C1 => n180, C2 => 
                           MEM_IN(27), A => n9310, ZN => n9309);
   U10341 : OAI22_X1 port map( A1 => n10898, A2 => n281, B1 => n5141, B2 => 
                           n133, ZN => n9310);
   U10342 : AOI22_X1 port map( A1 => n9199, A2 => n5142, B1 => n9200, B2 => 
                           n5143, ZN => n9308);
   U10343 : AOI22_X1 port map( A1 => n9201, A2 => n5144, B1 => n9202, B2 => 
                           n5145, ZN => n9307);
   U10344 : NAND3_X1 port map( A1 => n9311, A2 => n9312, A3 => n9313, ZN => 
                           n12260_port);
   U10345 : AOI221_X1 port map( B1 => n9196, B2 => n5149, C1 => n180, C2 => 
                           MEM_IN(28), A => n9314, ZN => n9313);
   U10346 : OAI22_X1 port map( A1 => n10897, A2 => n281, B1 => n5151, B2 => 
                           n133, ZN => n9314);
   U10347 : AOI22_X1 port map( A1 => n9199, A2 => n5152, B1 => n9200, B2 => 
                           n5153, ZN => n9312);
   U10348 : AOI22_X1 port map( A1 => n9201, A2 => n5154, B1 => n9202, B2 => 
                           n5155, ZN => n9311);
   U10349 : NAND3_X1 port map( A1 => n9315, A2 => n9316, A3 => n9317, ZN => 
                           n12259_port);
   U10350 : AOI221_X1 port map( B1 => n9196, B2 => n5159, C1 => n180, C2 => 
                           MEM_IN(29), A => n9318, ZN => n9317);
   U10351 : OAI22_X1 port map( A1 => n10896, A2 => n281, B1 => n5161, B2 => 
                           n133, ZN => n9318);
   U10352 : AOI22_X1 port map( A1 => n9199, A2 => n5162, B1 => n9200, B2 => 
                           n5163, ZN => n9316);
   U10353 : AOI22_X1 port map( A1 => n9201, A2 => n5164, B1 => n9202, B2 => 
                           n5165, ZN => n9315);
   U10354 : NAND3_X1 port map( A1 => n9319, A2 => n9320, A3 => n9321, ZN => 
                           n12258_port);
   U10355 : AOI221_X1 port map( B1 => n9196, B2 => n5169, C1 => n180, C2 => 
                           MEM_IN(30), A => n9322, ZN => n9321);
   U10356 : OAI22_X1 port map( A1 => n10895, A2 => n281, B1 => n5171, B2 => 
                           n133, ZN => n9322);
   U10357 : AOI22_X1 port map( A1 => n9199, A2 => n5172, B1 => n9200, B2 => 
                           n5173, ZN => n9320);
   U10358 : AOI22_X1 port map( A1 => n9201, A2 => n5174, B1 => n9202, B2 => 
                           n5175, ZN => n9319);
   U10359 : NAND3_X1 port map( A1 => n9323, A2 => n9324, A3 => n9325, ZN => 
                           n12257_port);
   U10360 : AOI221_X1 port map( B1 => n9196, B2 => n5179, C1 => n180, C2 => 
                           MEM_IN(31), A => n9326, ZN => n9325);
   U10361 : OAI22_X1 port map( A1 => n10894, A2 => n281, B1 => n5181, B2 => 
                           n133, ZN => n9326);
   U10362 : INV_X1 port map( A => n9330, ZN => n9329);
   U10363 : NAND2_X1 port map( A1 => n5206, A2 => n9036, ZN => n9031);
   U10364 : NAND2_X1 port map( A1 => n8740, A2 => n5206, ZN => n9036);
   U10365 : AOI22_X1 port map( A1 => n9199, A2 => n5191, B1 => n9200, B2 => 
                           n5192, ZN => n9324);
   U10366 : AOI22_X1 port map( A1 => n9201, A2 => n5195, B1 => n9202, B2 => 
                           n5196, ZN => n9323);
   U10367 : OAI22_X1 port map( A1 => n9330, A2 => n9328, B1 => n208, B2 => n280
                           , ZN => n9331);
   U10368 : NAND3_X1 port map( A1 => n208, A2 => n281, A3 => n8302, ZN => n9328
                           );
   U10369 : INV_X1 port map( A => n9327, ZN => n8302);
   U10370 : OAI22_X1 port map( A1 => n4786, A2 => n9334, B1 => n9335, B2 => 
                           n5204, ZN => n9198);
   U10371 : NOR2_X1 port map( A1 => n9327, A2 => n9330, ZN => n9335);
   U10372 : NAND2_X1 port map( A1 => n9336, A2 => n8889, ZN => n9327);
   U10373 : AOI211_X1 port map( C1 => n8891, C2 => n9337, A => n9190, B => 
                           n9333, ZN => n9334);
   U10374 : OAI21_X1 port map( B1 => n8889, B2 => n4787, A => n5368, ZN => 
                           n9190);
   U10375 : AND2_X1 port map( A1 => n8740, A2 => n8745, ZN => n8889);
   U10376 : AND2_X1 port map( A1 => n8596, A2 => n8450, ZN => n8740);
   U10377 : INV_X1 port map( A => n9043, ZN => n8891);
   U10378 : NAND2_X1 port map( A1 => n9338, A2 => n9339, ZN => n9330);
   U10379 : NOR2_X1 port map( A1 => n8450, A2 => n4787, ZN => n8886);
   U10380 : NAND2_X1 port map( A1 => n8895, A2 => n5775, ZN => n8450);
   U10381 : NAND3_X1 port map( A1 => n9340, A2 => n9341, A3 => n9342, ZN => 
                           n12256_port);
   U10382 : AOI221_X1 port map( B1 => n212, B2 => n4863, C1 => n181, C2 => 
                           MEM_IN(0), A => n9343, ZN => n9342);
   U10383 : OAI22_X1 port map( A1 => n10893, A2 => n255, B1 => n4867, B2 => 
                           n130, ZN => n9343);
   U10384 : AOI22_X1 port map( A1 => n195, A2 => n4869, B1 => n157, B2 => n4871
                           , ZN => n9341);
   U10385 : AOI22_X1 port map( A1 => n237, A2 => n4873, B1 => n154, B2 => n4875
                           , ZN => n9340);
   U10386 : NAND3_X1 port map( A1 => n9345, A2 => n9346, A3 => n9347, ZN => 
                           n12255_port);
   U10387 : AOI221_X1 port map( B1 => n212, B2 => n4879, C1 => n181, C2 => 
                           MEM_IN(1), A => n9348, ZN => n9347);
   U10388 : OAI22_X1 port map( A1 => n10892, A2 => n255, B1 => n4881, B2 => 
                           n130, ZN => n9348);
   U10389 : AOI22_X1 port map( A1 => n195, A2 => n4882, B1 => n157, B2 => n4883
                           , ZN => n9346);
   U10390 : AOI22_X1 port map( A1 => n237, A2 => n4884, B1 => n154, B2 => n4885
                           , ZN => n9345);
   U10391 : NAND3_X1 port map( A1 => n9349, A2 => n9350, A3 => n9351, ZN => 
                           n12254_port);
   U10392 : AOI221_X1 port map( B1 => n212, B2 => n4889, C1 => n181, C2 => 
                           MEM_IN(2), A => n9352, ZN => n9351);
   U10393 : OAI22_X1 port map( A1 => n10891, A2 => n255, B1 => n4891, B2 => 
                           n130, ZN => n9352);
   U10394 : AOI22_X1 port map( A1 => n195, A2 => n4892, B1 => n157, B2 => n4893
                           , ZN => n9350);
   U10395 : AOI22_X1 port map( A1 => n237, A2 => n4894, B1 => n154, B2 => n4895
                           , ZN => n9349);
   U10396 : NAND3_X1 port map( A1 => n9353, A2 => n9354, A3 => n9355, ZN => 
                           n12253_port);
   U10397 : AOI221_X1 port map( B1 => n212, B2 => n4899, C1 => n181, C2 => 
                           MEM_IN(3), A => n9356, ZN => n9355);
   U10398 : OAI22_X1 port map( A1 => n10890, A2 => n255, B1 => n4901, B2 => 
                           n130, ZN => n9356);
   U10399 : AOI22_X1 port map( A1 => n195, A2 => n4902, B1 => n157, B2 => n4903
                           , ZN => n9354);
   U10400 : AOI22_X1 port map( A1 => n237, A2 => n4904, B1 => n154, B2 => n4905
                           , ZN => n9353);
   U10401 : NAND3_X1 port map( A1 => n9357, A2 => n9358, A3 => n9359, ZN => 
                           n12252_port);
   U10402 : AOI221_X1 port map( B1 => n212, B2 => n4909, C1 => n181, C2 => 
                           MEM_IN(4), A => n9360, ZN => n9359);
   U10403 : OAI22_X1 port map( A1 => n10889, A2 => n255, B1 => n4911, B2 => 
                           n130, ZN => n9360);
   U10404 : AOI22_X1 port map( A1 => n195, A2 => n4912, B1 => n157, B2 => n4913
                           , ZN => n9358);
   U10405 : AOI22_X1 port map( A1 => n237, A2 => n4914, B1 => n154, B2 => n4915
                           , ZN => n9357);
   U10406 : NAND3_X1 port map( A1 => n9361, A2 => n9362, A3 => n9363, ZN => 
                           n12251_port);
   U10407 : AOI221_X1 port map( B1 => n212, B2 => n4919, C1 => n181, C2 => 
                           MEM_IN(5), A => n9364, ZN => n9363);
   U10408 : OAI22_X1 port map( A1 => n10888, A2 => n255, B1 => n4921, B2 => 
                           n130, ZN => n9364);
   U10409 : AOI22_X1 port map( A1 => n195, A2 => n4922, B1 => n157, B2 => n4923
                           , ZN => n9362);
   U10410 : AOI22_X1 port map( A1 => n237, A2 => n4924, B1 => n154, B2 => n4925
                           , ZN => n9361);
   U10411 : NAND3_X1 port map( A1 => n9365, A2 => n9366, A3 => n9367, ZN => 
                           n12250_port);
   U10412 : AOI221_X1 port map( B1 => n212, B2 => n4929, C1 => n181, C2 => 
                           MEM_IN(6), A => n9368, ZN => n9367);
   U10413 : OAI22_X1 port map( A1 => n10887, A2 => n255, B1 => n4931, B2 => 
                           n130, ZN => n9368);
   U10414 : AOI22_X1 port map( A1 => n195, A2 => n4932, B1 => n157, B2 => n4933
                           , ZN => n9366);
   U10415 : AOI22_X1 port map( A1 => n237, A2 => n4934, B1 => n154, B2 => n4935
                           , ZN => n9365);
   U10416 : NAND3_X1 port map( A1 => n9369, A2 => n9370, A3 => n9371, ZN => 
                           n12249_port);
   U10417 : AOI221_X1 port map( B1 => n212, B2 => n4939, C1 => n181, C2 => 
                           MEM_IN(7), A => n9372, ZN => n9371);
   U10418 : OAI22_X1 port map( A1 => n10886, A2 => n255, B1 => n4941, B2 => 
                           n130, ZN => n9372);
   U10419 : AOI22_X1 port map( A1 => n195, A2 => n4942, B1 => n157, B2 => n4943
                           , ZN => n9370);
   U10420 : AOI22_X1 port map( A1 => n237, A2 => n4944, B1 => n154, B2 => n4945
                           , ZN => n9369);
   U10421 : NAND3_X1 port map( A1 => n9373, A2 => n9374, A3 => n9375, ZN => 
                           n12248_port);
   U10422 : AOI221_X1 port map( B1 => n212, B2 => n4949, C1 => n181, C2 => 
                           MEM_IN(8), A => n9376, ZN => n9375);
   U10423 : OAI22_X1 port map( A1 => n10885, A2 => n255, B1 => n4951, B2 => 
                           n130, ZN => n9376);
   U10424 : AOI22_X1 port map( A1 => n195, A2 => n4952, B1 => n157, B2 => n4953
                           , ZN => n9374);
   U10425 : AOI22_X1 port map( A1 => n237, A2 => n4954, B1 => n154, B2 => n4955
                           , ZN => n9373);
   U10426 : NAND3_X1 port map( A1 => n9377, A2 => n9378, A3 => n9379, ZN => 
                           n12247_port);
   U10427 : AOI221_X1 port map( B1 => n212, B2 => n4959, C1 => n181, C2 => 
                           MEM_IN(9), A => n9380, ZN => n9379);
   U10428 : OAI22_X1 port map( A1 => n10884, A2 => n255, B1 => n4961, B2 => 
                           n130, ZN => n9380);
   U10429 : AOI22_X1 port map( A1 => n195, A2 => n4962, B1 => n157, B2 => n4963
                           , ZN => n9378);
   U10430 : AOI22_X1 port map( A1 => n237, A2 => n4964, B1 => n154, B2 => n4965
                           , ZN => n9377);
   U10431 : NAND3_X1 port map( A1 => n9381, A2 => n9382, A3 => n9383, ZN => 
                           n12246_port);
   U10432 : AOI221_X1 port map( B1 => n212, B2 => n4969, C1 => n181, C2 => 
                           MEM_IN(10), A => n9384, ZN => n9383);
   U10433 : OAI22_X1 port map( A1 => n10883, A2 => n255, B1 => n4971, B2 => 
                           n130, ZN => n9384);
   U10434 : AOI22_X1 port map( A1 => n195, A2 => n4972, B1 => n157, B2 => n4973
                           , ZN => n9382);
   U10435 : AOI22_X1 port map( A1 => n237, A2 => n4974, B1 => n154, B2 => n4975
                           , ZN => n9381);
   U10436 : NAND3_X1 port map( A1 => n9385, A2 => n9386, A3 => n9387, ZN => 
                           n12245_port);
   U10437 : AOI221_X1 port map( B1 => n212, B2 => n4979, C1 => n181, C2 => 
                           MEM_IN(11), A => n9388, ZN => n9387);
   U10438 : OAI22_X1 port map( A1 => n10882, A2 => n255, B1 => n4981, B2 => 
                           n130, ZN => n9388);
   U10439 : AOI22_X1 port map( A1 => n195, A2 => n4982, B1 => n157, B2 => n4983
                           , ZN => n9386);
   U10440 : AOI22_X1 port map( A1 => n237, A2 => n4984, B1 => n154, B2 => n4985
                           , ZN => n9385);
   U10441 : NAND3_X1 port map( A1 => n9389, A2 => n9390, A3 => n9391, ZN => 
                           n12244_port);
   U10442 : AOI221_X1 port map( B1 => n212, B2 => n4989, C1 => n181, C2 => 
                           MEM_IN(12), A => n9392, ZN => n9391);
   U10443 : OAI22_X1 port map( A1 => n10881, A2 => n255, B1 => n4991, B2 => 
                           n130, ZN => n9392);
   U10444 : AOI22_X1 port map( A1 => n195, A2 => n4992, B1 => n157, B2 => n4993
                           , ZN => n9390);
   U10445 : AOI22_X1 port map( A1 => n237, A2 => n4994, B1 => n154, B2 => n4995
                           , ZN => n9389);
   U10446 : NAND3_X1 port map( A1 => n9393, A2 => n9394, A3 => n9395, ZN => 
                           n12243_port);
   U10447 : AOI221_X1 port map( B1 => n212, B2 => n4999, C1 => n181, C2 => 
                           MEM_IN(13), A => n9396, ZN => n9395);
   U10448 : OAI22_X1 port map( A1 => n10880, A2 => n255, B1 => n5001, B2 => 
                           n130, ZN => n9396);
   U10449 : AOI22_X1 port map( A1 => n195, A2 => n5002, B1 => n157, B2 => n5003
                           , ZN => n9394);
   U10450 : AOI22_X1 port map( A1 => n237, A2 => n5004, B1 => n154, B2 => n5005
                           , ZN => n9393);
   U10451 : NAND3_X1 port map( A1 => n9397, A2 => n9398, A3 => n9399, ZN => 
                           n12242_port);
   U10452 : AOI221_X1 port map( B1 => n212, B2 => n5009, C1 => n181, C2 => 
                           MEM_IN(14), A => n9400, ZN => n9399);
   U10453 : OAI22_X1 port map( A1 => n10879, A2 => n255, B1 => n5011, B2 => 
                           n130, ZN => n9400);
   U10454 : AOI22_X1 port map( A1 => n195, A2 => n5012, B1 => n157, B2 => n5013
                           , ZN => n9398);
   U10455 : AOI22_X1 port map( A1 => n237, A2 => n5014, B1 => n154, B2 => n5015
                           , ZN => n9397);
   U10456 : NAND3_X1 port map( A1 => n9401, A2 => n9402, A3 => n9403, ZN => 
                           n12241_port);
   U10457 : AOI221_X1 port map( B1 => n212, B2 => n5019, C1 => n181, C2 => 
                           MEM_IN(15), A => n9404, ZN => n9403);
   U10458 : OAI22_X1 port map( A1 => n10878, A2 => n255, B1 => n5021, B2 => 
                           n130, ZN => n9404);
   U10459 : AOI22_X1 port map( A1 => n195, A2 => n5022, B1 => n157, B2 => n5023
                           , ZN => n9402);
   U10460 : AOI22_X1 port map( A1 => n237, A2 => n5024, B1 => n154, B2 => n5025
                           , ZN => n9401);
   U10461 : NAND3_X1 port map( A1 => n9405, A2 => n9406, A3 => n9407, ZN => 
                           n12240_port);
   U10462 : AOI221_X1 port map( B1 => n212, B2 => n5029, C1 => n181, C2 => 
                           MEM_IN(16), A => n9408, ZN => n9407);
   U10463 : OAI22_X1 port map( A1 => n10877, A2 => n255, B1 => n5031, B2 => 
                           n130, ZN => n9408);
   U10464 : AOI22_X1 port map( A1 => n195, A2 => n5032, B1 => n157, B2 => n5033
                           , ZN => n9406);
   U10465 : AOI22_X1 port map( A1 => n237, A2 => n5034, B1 => n154, B2 => n5035
                           , ZN => n9405);
   U10466 : NAND3_X1 port map( A1 => n9409, A2 => n9410, A3 => n9411, ZN => 
                           n12239_port);
   U10467 : AOI221_X1 port map( B1 => n212, B2 => n5039, C1 => n181, C2 => 
                           MEM_IN(17), A => n9412, ZN => n9411);
   U10468 : OAI22_X1 port map( A1 => n10876, A2 => n255, B1 => n5041, B2 => 
                           n130, ZN => n9412);
   U10469 : AOI22_X1 port map( A1 => n195, A2 => n5042, B1 => n157, B2 => n5043
                           , ZN => n9410);
   U10470 : AOI22_X1 port map( A1 => n237, A2 => n5044, B1 => n154, B2 => n5045
                           , ZN => n9409);
   U10471 : NAND3_X1 port map( A1 => n9413, A2 => n9414, A3 => n9415, ZN => 
                           n12238_port);
   U10472 : AOI221_X1 port map( B1 => n212, B2 => n5049, C1 => n181, C2 => 
                           MEM_IN(18), A => n9416, ZN => n9415);
   U10473 : OAI22_X1 port map( A1 => n10875, A2 => n255, B1 => n5051, B2 => 
                           n130, ZN => n9416);
   U10474 : AOI22_X1 port map( A1 => n195, A2 => n5052, B1 => n157, B2 => n5053
                           , ZN => n9414);
   U10475 : AOI22_X1 port map( A1 => n237, A2 => n5054, B1 => n154, B2 => n5055
                           , ZN => n9413);
   U10476 : NAND3_X1 port map( A1 => n9417, A2 => n9418, A3 => n9419, ZN => 
                           n12237_port);
   U10477 : AOI221_X1 port map( B1 => n212, B2 => n5059, C1 => n181, C2 => 
                           MEM_IN(19), A => n9420, ZN => n9419);
   U10478 : OAI22_X1 port map( A1 => n10874, A2 => n255, B1 => n5061, B2 => 
                           n130, ZN => n9420);
   U10479 : AOI22_X1 port map( A1 => n195, A2 => n5062, B1 => n157, B2 => n5063
                           , ZN => n9418);
   U10480 : AOI22_X1 port map( A1 => n237, A2 => n5064, B1 => n154, B2 => n5065
                           , ZN => n9417);
   U10481 : NAND3_X1 port map( A1 => n9421, A2 => n9422, A3 => n9423, ZN => 
                           n12236_port);
   U10482 : AOI221_X1 port map( B1 => n212, B2 => n5069, C1 => n181, C2 => 
                           MEM_IN(20), A => n9424, ZN => n9423);
   U10483 : OAI22_X1 port map( A1 => n10873, A2 => n255, B1 => n5071, B2 => 
                           n130, ZN => n9424);
   U10484 : AOI22_X1 port map( A1 => n195, A2 => n5072, B1 => n157, B2 => n5073
                           , ZN => n9422);
   U10485 : AOI22_X1 port map( A1 => n237, A2 => n5074, B1 => n154, B2 => n5075
                           , ZN => n9421);
   U10486 : NAND3_X1 port map( A1 => n9425, A2 => n9426, A3 => n9427, ZN => 
                           n12235_port);
   U10487 : AOI221_X1 port map( B1 => n212, B2 => n5079, C1 => n181, C2 => 
                           MEM_IN(21), A => n9428, ZN => n9427);
   U10488 : OAI22_X1 port map( A1 => n10872, A2 => n255, B1 => n5081, B2 => 
                           n130, ZN => n9428);
   U10489 : AOI22_X1 port map( A1 => n195, A2 => n5082, B1 => n157, B2 => n5083
                           , ZN => n9426);
   U10490 : AOI22_X1 port map( A1 => n237, A2 => n5084, B1 => n154, B2 => n5085
                           , ZN => n9425);
   U10491 : NAND3_X1 port map( A1 => n9429, A2 => n9430, A3 => n9431, ZN => 
                           n12234_port);
   U10492 : AOI221_X1 port map( B1 => n212, B2 => n5089, C1 => n181, C2 => 
                           MEM_IN(22), A => n9432, ZN => n9431);
   U10493 : OAI22_X1 port map( A1 => n10871, A2 => n255, B1 => n5091, B2 => 
                           n130, ZN => n9432);
   U10494 : AOI22_X1 port map( A1 => n195, A2 => n5092, B1 => n157, B2 => n5093
                           , ZN => n9430);
   U10495 : AOI22_X1 port map( A1 => n237, A2 => n5094, B1 => n154, B2 => n5095
                           , ZN => n9429);
   U10496 : NAND3_X1 port map( A1 => n9433, A2 => n9434, A3 => n9435, ZN => 
                           n12233_port);
   U10497 : AOI221_X1 port map( B1 => n212, B2 => n5099, C1 => n181, C2 => 
                           MEM_IN(23), A => n9436, ZN => n9435);
   U10498 : OAI22_X1 port map( A1 => n10870, A2 => n255, B1 => n5101, B2 => 
                           n130, ZN => n9436);
   U10499 : AOI22_X1 port map( A1 => n195, A2 => n5102, B1 => n157, B2 => n5103
                           , ZN => n9434);
   U10500 : AOI22_X1 port map( A1 => n237, A2 => n5104, B1 => n154, B2 => n5105
                           , ZN => n9433);
   U10501 : NAND3_X1 port map( A1 => n9437, A2 => n9438, A3 => n9439, ZN => 
                           n12232_port);
   U10502 : AOI221_X1 port map( B1 => n212, B2 => n5109, C1 => n181, C2 => 
                           MEM_IN(24), A => n9440, ZN => n9439);
   U10503 : OAI22_X1 port map( A1 => n10869, A2 => n255, B1 => n5111, B2 => 
                           n130, ZN => n9440);
   U10504 : AOI22_X1 port map( A1 => n195, A2 => n5112, B1 => n157, B2 => n5113
                           , ZN => n9438);
   U10505 : AOI22_X1 port map( A1 => n237, A2 => n5114, B1 => n154, B2 => n5115
                           , ZN => n9437);
   U10506 : NAND3_X1 port map( A1 => n9441, A2 => n9442, A3 => n9443, ZN => 
                           n12231_port);
   U10507 : AOI221_X1 port map( B1 => n212, B2 => n5119, C1 => n181, C2 => 
                           MEM_IN(25), A => n9444, ZN => n9443);
   U10508 : OAI22_X1 port map( A1 => n10868, A2 => n255, B1 => n5121, B2 => 
                           n130, ZN => n9444);
   U10509 : AOI22_X1 port map( A1 => n195, A2 => n5122, B1 => n157, B2 => n5123
                           , ZN => n9442);
   U10510 : AOI22_X1 port map( A1 => n237, A2 => n5124, B1 => n154, B2 => n5125
                           , ZN => n9441);
   U10511 : NAND3_X1 port map( A1 => n9445, A2 => n9446, A3 => n9447, ZN => 
                           n12230_port);
   U10512 : AOI221_X1 port map( B1 => n212, B2 => n5129, C1 => n181, C2 => 
                           MEM_IN(26), A => n9448, ZN => n9447);
   U10513 : OAI22_X1 port map( A1 => n10867, A2 => n255, B1 => n5131, B2 => 
                           n130, ZN => n9448);
   U10514 : AOI22_X1 port map( A1 => n195, A2 => n5132, B1 => n157, B2 => n5133
                           , ZN => n9446);
   U10515 : AOI22_X1 port map( A1 => n237, A2 => n5134, B1 => n154, B2 => n5135
                           , ZN => n9445);
   U10516 : NAND3_X1 port map( A1 => n9449, A2 => n9450, A3 => n9451, ZN => 
                           n12229_port);
   U10517 : AOI221_X1 port map( B1 => n212, B2 => n5139, C1 => n181, C2 => 
                           MEM_IN(27), A => n9452, ZN => n9451);
   U10518 : OAI22_X1 port map( A1 => n10866, A2 => n255, B1 => n5141, B2 => 
                           n130, ZN => n9452);
   U10519 : AOI22_X1 port map( A1 => n195, A2 => n5142, B1 => n157, B2 => n5143
                           , ZN => n9450);
   U10520 : AOI22_X1 port map( A1 => n237, A2 => n5144, B1 => n154, B2 => n5145
                           , ZN => n9449);
   U10521 : NAND3_X1 port map( A1 => n9453, A2 => n9454, A3 => n9455, ZN => 
                           n12228_port);
   U10522 : AOI221_X1 port map( B1 => n212, B2 => n5149, C1 => n181, C2 => 
                           MEM_IN(28), A => n9456, ZN => n9455);
   U10523 : OAI22_X1 port map( A1 => n10865, A2 => n255, B1 => n5151, B2 => 
                           n130, ZN => n9456);
   U10524 : AOI22_X1 port map( A1 => n195, A2 => n5152, B1 => n157, B2 => n5153
                           , ZN => n9454);
   U10525 : AOI22_X1 port map( A1 => n237, A2 => n5154, B1 => n154, B2 => n5155
                           , ZN => n9453);
   U10526 : NAND3_X1 port map( A1 => n9457, A2 => n9458, A3 => n9459, ZN => 
                           n12227_port);
   U10527 : AOI221_X1 port map( B1 => n212, B2 => n5159, C1 => n181, C2 => 
                           MEM_IN(29), A => n9460, ZN => n9459);
   U10528 : OAI22_X1 port map( A1 => n10864, A2 => n255, B1 => n5161, B2 => 
                           n130, ZN => n9460);
   U10529 : AOI22_X1 port map( A1 => n195, A2 => n5162, B1 => n157, B2 => n5163
                           , ZN => n9458);
   U10530 : AOI22_X1 port map( A1 => n237, A2 => n5164, B1 => n154, B2 => n5165
                           , ZN => n9457);
   U10531 : NAND3_X1 port map( A1 => n9461, A2 => n9462, A3 => n9463, ZN => 
                           n12226_port);
   U10532 : AOI221_X1 port map( B1 => n212, B2 => n5169, C1 => n181, C2 => 
                           MEM_IN(30), A => n9464, ZN => n9463);
   U10533 : OAI22_X1 port map( A1 => n10863, A2 => n255, B1 => n5171, B2 => 
                           n130, ZN => n9464);
   U10534 : AOI22_X1 port map( A1 => n195, A2 => n5172, B1 => n157, B2 => n5173
                           , ZN => n9462);
   U10535 : AOI22_X1 port map( A1 => n237, A2 => n5174, B1 => n154, B2 => n5175
                           , ZN => n9461);
   U10536 : NAND3_X1 port map( A1 => n9465, A2 => n9466, A3 => n9467, ZN => 
                           n12225_port);
   U10537 : AOI221_X1 port map( B1 => n212, B2 => n5179, C1 => n181, C2 => 
                           MEM_IN(31), A => n9468, ZN => n9467);
   U10538 : OAI22_X1 port map( A1 => n10862, A2 => n255, B1 => n5181, B2 => 
                           n130, ZN => n9468);
   U10539 : INV_X1 port map( A => n9474, ZN => n9473);
   U10540 : AOI22_X1 port map( A1 => n195, A2 => n5191, B1 => n157, B2 => n5192
                           , ZN => n9466);
   U10541 : INV_X1 port map( A => n9333, ZN => n9332);
   U10542 : AOI22_X1 port map( A1 => n237, A2 => n5195, B1 => n154, B2 => n5196
                           , ZN => n9465);
   U10543 : AOI22_X1 port map( A1 => n9471, A2 => n9477, B1 => n4841, B2 => 
                           n255, ZN => n9472);
   U10544 : INV_X1 port map( A => n9470, ZN => n9477);
   U10545 : NAND3_X1 port map( A1 => n208, A2 => n255, A3 => n8449, ZN => n9470
                           );
   U10546 : INV_X1 port map( A => n9469, ZN => n8449);
   U10547 : OAI22_X1 port map( A1 => n4786, A2 => n9478, B1 => n9479, B2 => 
                           n5204, ZN => n9344);
   U10548 : NOR2_X1 port map( A1 => n9469, A2 => n9480, ZN => n9479);
   U10549 : NAND4_X1 port map( A1 => n9336, A2 => n9339, A3 => n8745, A4 => 
                           n8596, ZN => n9469);
   U10550 : NOR4_X1 port map( A1 => n9481, A2 => n9333, A3 => RESET, A4 => 
                           n9482, ZN => n9478);
   U10551 : OAI211_X1 port map( C1 => n5923, C2 => n9043, A => n9033, B => 
                           n9185, ZN => n9481);
   U10552 : INV_X1 port map( A => n9186, ZN => n9185);
   U10553 : INV_X1 port map( A => n9042, ZN => n9033);
   U10554 : NOR2_X1 port map( A1 => n8596, A2 => n4787, ZN => n9042);
   U10555 : INV_X1 port map( A => n9480, ZN => n9471);
   U10556 : NAND2_X1 port map( A1 => n9483, A2 => n9484, ZN => n9480);
   U10557 : NAND2_X1 port map( A1 => n8895, A2 => n5926, ZN => n8596);
   U10558 : NAND3_X1 port map( A1 => n9485, A2 => n9486, A3 => n9487, ZN => 
                           n12224_port);
   U10559 : AOI221_X1 port map( B1 => n9488, B2 => n4863, C1 => n176, C2 => 
                           MEM_IN(0), A => n9489, ZN => n9487);
   U10560 : OAI22_X1 port map( A1 => n10861, A2 => n283, B1 => n4867, B2 => 
                           n131, ZN => n9489);
   U10561 : AOI22_X1 port map( A1 => n9491, A2 => n4869, B1 => n9492, B2 => 
                           n4871, ZN => n9486);
   U10562 : AOI22_X1 port map( A1 => n9493, A2 => n4873, B1 => n9494, B2 => 
                           n4875, ZN => n9485);
   U10563 : NAND3_X1 port map( A1 => n9495, A2 => n9496, A3 => n9497, ZN => 
                           n12223_port);
   U10564 : AOI221_X1 port map( B1 => n9488, B2 => n4879, C1 => n176, C2 => 
                           MEM_IN(1), A => n9498, ZN => n9497);
   U10565 : OAI22_X1 port map( A1 => n10860, A2 => n283, B1 => n4881, B2 => 
                           n131, ZN => n9498);
   U10566 : AOI22_X1 port map( A1 => n9491, A2 => n4882, B1 => n9492, B2 => 
                           n4883, ZN => n9496);
   U10567 : AOI22_X1 port map( A1 => n9493, A2 => n4884, B1 => n9494, B2 => 
                           n4885, ZN => n9495);
   U10568 : NAND3_X1 port map( A1 => n9499, A2 => n9500, A3 => n9501, ZN => 
                           n12222_port);
   U10569 : AOI221_X1 port map( B1 => n9488, B2 => n4889, C1 => n176, C2 => 
                           MEM_IN(2), A => n9502, ZN => n9501);
   U10570 : OAI22_X1 port map( A1 => n10859, A2 => n283, B1 => n4891, B2 => 
                           n131, ZN => n9502);
   U10571 : AOI22_X1 port map( A1 => n9491, A2 => n4892, B1 => n9492, B2 => 
                           n4893, ZN => n9500);
   U10572 : AOI22_X1 port map( A1 => n9493, A2 => n4894, B1 => n9494, B2 => 
                           n4895, ZN => n9499);
   U10573 : NAND3_X1 port map( A1 => n9503, A2 => n9504, A3 => n9505, ZN => 
                           n12221_port);
   U10574 : AOI221_X1 port map( B1 => n9488, B2 => n4899, C1 => n176, C2 => 
                           MEM_IN(3), A => n9506, ZN => n9505);
   U10575 : OAI22_X1 port map( A1 => n10858, A2 => n283, B1 => n4901, B2 => 
                           n131, ZN => n9506);
   U10576 : AOI22_X1 port map( A1 => n9491, A2 => n4902, B1 => n9492, B2 => 
                           n4903, ZN => n9504);
   U10577 : AOI22_X1 port map( A1 => n9493, A2 => n4904, B1 => n9494, B2 => 
                           n4905, ZN => n9503);
   U10578 : NAND3_X1 port map( A1 => n9507, A2 => n9508, A3 => n9509, ZN => 
                           n12220_port);
   U10579 : AOI221_X1 port map( B1 => n9488, B2 => n4909, C1 => n176, C2 => 
                           MEM_IN(4), A => n9510, ZN => n9509);
   U10580 : OAI22_X1 port map( A1 => n10857, A2 => n283, B1 => n4911, B2 => 
                           n131, ZN => n9510);
   U10581 : AOI22_X1 port map( A1 => n9491, A2 => n4912, B1 => n9492, B2 => 
                           n4913, ZN => n9508);
   U10582 : AOI22_X1 port map( A1 => n9493, A2 => n4914, B1 => n9494, B2 => 
                           n4915, ZN => n9507);
   U10583 : NAND3_X1 port map( A1 => n9511, A2 => n9512, A3 => n9513, ZN => 
                           n12219_port);
   U10584 : AOI221_X1 port map( B1 => n9488, B2 => n4919, C1 => n176, C2 => 
                           MEM_IN(5), A => n9514, ZN => n9513);
   U10585 : OAI22_X1 port map( A1 => n10856, A2 => n283, B1 => n4921, B2 => 
                           n131, ZN => n9514);
   U10586 : AOI22_X1 port map( A1 => n9491, A2 => n4922, B1 => n9492, B2 => 
                           n4923, ZN => n9512);
   U10587 : AOI22_X1 port map( A1 => n9493, A2 => n4924, B1 => n9494, B2 => 
                           n4925, ZN => n9511);
   U10588 : NAND3_X1 port map( A1 => n9515, A2 => n9516, A3 => n9517, ZN => 
                           n12218_port);
   U10589 : AOI221_X1 port map( B1 => n9488, B2 => n4929, C1 => n176, C2 => 
                           MEM_IN(6), A => n9518, ZN => n9517);
   U10590 : OAI22_X1 port map( A1 => n10855, A2 => n283, B1 => n4931, B2 => 
                           n131, ZN => n9518);
   U10591 : AOI22_X1 port map( A1 => n9491, A2 => n4932, B1 => n9492, B2 => 
                           n4933, ZN => n9516);
   U10592 : AOI22_X1 port map( A1 => n9493, A2 => n4934, B1 => n9494, B2 => 
                           n4935, ZN => n9515);
   U10593 : NAND3_X1 port map( A1 => n9519, A2 => n9520, A3 => n9521, ZN => 
                           n12217_port);
   U10594 : AOI221_X1 port map( B1 => n9488, B2 => n4939, C1 => n176, C2 => 
                           MEM_IN(7), A => n9522, ZN => n9521);
   U10595 : OAI22_X1 port map( A1 => n10854, A2 => n283, B1 => n4941, B2 => 
                           n131, ZN => n9522);
   U10596 : AOI22_X1 port map( A1 => n9491, A2 => n4942, B1 => n9492, B2 => 
                           n4943, ZN => n9520);
   U10597 : AOI22_X1 port map( A1 => n9493, A2 => n4944, B1 => n9494, B2 => 
                           n4945, ZN => n9519);
   U10598 : NAND3_X1 port map( A1 => n9523, A2 => n9524, A3 => n9525, ZN => 
                           n12216_port);
   U10599 : AOI221_X1 port map( B1 => n9488, B2 => n4949, C1 => n176, C2 => 
                           MEM_IN(8), A => n9526, ZN => n9525);
   U10600 : OAI22_X1 port map( A1 => n10853, A2 => n283, B1 => n4951, B2 => 
                           n131, ZN => n9526);
   U10601 : AOI22_X1 port map( A1 => n9491, A2 => n4952, B1 => n9492, B2 => 
                           n4953, ZN => n9524);
   U10602 : AOI22_X1 port map( A1 => n9493, A2 => n4954, B1 => n9494, B2 => 
                           n4955, ZN => n9523);
   U10603 : NAND3_X1 port map( A1 => n9527, A2 => n9528, A3 => n9529, ZN => 
                           n12215_port);
   U10604 : AOI221_X1 port map( B1 => n9488, B2 => n4959, C1 => n176, C2 => 
                           MEM_IN(9), A => n9530, ZN => n9529);
   U10605 : OAI22_X1 port map( A1 => n10852, A2 => n283, B1 => n4961, B2 => 
                           n131, ZN => n9530);
   U10606 : AOI22_X1 port map( A1 => n9491, A2 => n4962, B1 => n9492, B2 => 
                           n4963, ZN => n9528);
   U10607 : AOI22_X1 port map( A1 => n9493, A2 => n4964, B1 => n9494, B2 => 
                           n4965, ZN => n9527);
   U10608 : NAND3_X1 port map( A1 => n9531, A2 => n9532, A3 => n9533, ZN => 
                           n12214_port);
   U10609 : AOI221_X1 port map( B1 => n9488, B2 => n4969, C1 => n176, C2 => 
                           MEM_IN(10), A => n9534, ZN => n9533);
   U10610 : OAI22_X1 port map( A1 => n10851, A2 => n283, B1 => n4971, B2 => 
                           n131, ZN => n9534);
   U10611 : AOI22_X1 port map( A1 => n9491, A2 => n4972, B1 => n9492, B2 => 
                           n4973, ZN => n9532);
   U10612 : AOI22_X1 port map( A1 => n9493, A2 => n4974, B1 => n9494, B2 => 
                           n4975, ZN => n9531);
   U10613 : NAND3_X1 port map( A1 => n9535, A2 => n9536, A3 => n9537, ZN => 
                           n12213_port);
   U10614 : AOI221_X1 port map( B1 => n9488, B2 => n4979, C1 => n176, C2 => 
                           MEM_IN(11), A => n9538, ZN => n9537);
   U10615 : OAI22_X1 port map( A1 => n10850, A2 => n283, B1 => n4981, B2 => 
                           n131, ZN => n9538);
   U10616 : AOI22_X1 port map( A1 => n9491, A2 => n4982, B1 => n9492, B2 => 
                           n4983, ZN => n9536);
   U10617 : AOI22_X1 port map( A1 => n9493, A2 => n4984, B1 => n9494, B2 => 
                           n4985, ZN => n9535);
   U10618 : NAND3_X1 port map( A1 => n9539, A2 => n9540, A3 => n9541, ZN => 
                           n12212_port);
   U10619 : AOI221_X1 port map( B1 => n9488, B2 => n4989, C1 => n176, C2 => 
                           MEM_IN(12), A => n9542, ZN => n9541);
   U10620 : OAI22_X1 port map( A1 => n10849, A2 => n283, B1 => n4991, B2 => 
                           n131, ZN => n9542);
   U10621 : AOI22_X1 port map( A1 => n9491, A2 => n4992, B1 => n9492, B2 => 
                           n4993, ZN => n9540);
   U10622 : AOI22_X1 port map( A1 => n9493, A2 => n4994, B1 => n9494, B2 => 
                           n4995, ZN => n9539);
   U10623 : NAND3_X1 port map( A1 => n9543, A2 => n9544, A3 => n9545, ZN => 
                           n12211_port);
   U10624 : AOI221_X1 port map( B1 => n9488, B2 => n4999, C1 => n176, C2 => 
                           MEM_IN(13), A => n9546, ZN => n9545);
   U10625 : OAI22_X1 port map( A1 => n10848, A2 => n283, B1 => n5001, B2 => 
                           n131, ZN => n9546);
   U10626 : AOI22_X1 port map( A1 => n9491, A2 => n5002, B1 => n9492, B2 => 
                           n5003, ZN => n9544);
   U10627 : AOI22_X1 port map( A1 => n9493, A2 => n5004, B1 => n9494, B2 => 
                           n5005, ZN => n9543);
   U10628 : NAND3_X1 port map( A1 => n9547, A2 => n9548, A3 => n9549, ZN => 
                           n12210_port);
   U10629 : AOI221_X1 port map( B1 => n9488, B2 => n5009, C1 => n176, C2 => 
                           MEM_IN(14), A => n9550, ZN => n9549);
   U10630 : OAI22_X1 port map( A1 => n10847, A2 => n283, B1 => n5011, B2 => 
                           n131, ZN => n9550);
   U10631 : AOI22_X1 port map( A1 => n9491, A2 => n5012, B1 => n9492, B2 => 
                           n5013, ZN => n9548);
   U10632 : AOI22_X1 port map( A1 => n9493, A2 => n5014, B1 => n9494, B2 => 
                           n5015, ZN => n9547);
   U10633 : NAND3_X1 port map( A1 => n9551, A2 => n9552, A3 => n9553, ZN => 
                           n12209_port);
   U10634 : AOI221_X1 port map( B1 => n9488, B2 => n5019, C1 => n176, C2 => 
                           MEM_IN(15), A => n9554, ZN => n9553);
   U10635 : OAI22_X1 port map( A1 => n10846, A2 => n283, B1 => n5021, B2 => 
                           n131, ZN => n9554);
   U10636 : AOI22_X1 port map( A1 => n9491, A2 => n5022, B1 => n9492, B2 => 
                           n5023, ZN => n9552);
   U10637 : AOI22_X1 port map( A1 => n9493, A2 => n5024, B1 => n9494, B2 => 
                           n5025, ZN => n9551);
   U10638 : NAND3_X1 port map( A1 => n9555, A2 => n9556, A3 => n9557, ZN => 
                           n12208_port);
   U10639 : AOI221_X1 port map( B1 => n9488, B2 => n5029, C1 => n176, C2 => 
                           MEM_IN(16), A => n9558, ZN => n9557);
   U10640 : OAI22_X1 port map( A1 => n10845, A2 => n283, B1 => n5031, B2 => 
                           n131, ZN => n9558);
   U10641 : AOI22_X1 port map( A1 => n9491, A2 => n5032, B1 => n9492, B2 => 
                           n5033, ZN => n9556);
   U10642 : AOI22_X1 port map( A1 => n9493, A2 => n5034, B1 => n9494, B2 => 
                           n5035, ZN => n9555);
   U10643 : NAND3_X1 port map( A1 => n9559, A2 => n9560, A3 => n9561, ZN => 
                           n12207_port);
   U10644 : AOI221_X1 port map( B1 => n9488, B2 => n5039, C1 => n176, C2 => 
                           MEM_IN(17), A => n9562, ZN => n9561);
   U10645 : OAI22_X1 port map( A1 => n10844, A2 => n283, B1 => n5041, B2 => 
                           n131, ZN => n9562);
   U10646 : AOI22_X1 port map( A1 => n9491, A2 => n5042, B1 => n9492, B2 => 
                           n5043, ZN => n9560);
   U10647 : AOI22_X1 port map( A1 => n9493, A2 => n5044, B1 => n9494, B2 => 
                           n5045, ZN => n9559);
   U10648 : NAND3_X1 port map( A1 => n9563, A2 => n9564, A3 => n9565, ZN => 
                           n12206_port);
   U10649 : AOI221_X1 port map( B1 => n9488, B2 => n5049, C1 => n176, C2 => 
                           MEM_IN(18), A => n9566, ZN => n9565);
   U10650 : OAI22_X1 port map( A1 => n10843, A2 => n283, B1 => n5051, B2 => 
                           n131, ZN => n9566);
   U10651 : AOI22_X1 port map( A1 => n9491, A2 => n5052, B1 => n9492, B2 => 
                           n5053, ZN => n9564);
   U10652 : AOI22_X1 port map( A1 => n9493, A2 => n5054, B1 => n9494, B2 => 
                           n5055, ZN => n9563);
   U10653 : NAND3_X1 port map( A1 => n9567, A2 => n9568, A3 => n9569, ZN => 
                           n12205_port);
   U10654 : AOI221_X1 port map( B1 => n9488, B2 => n5059, C1 => n176, C2 => 
                           MEM_IN(19), A => n9570, ZN => n9569);
   U10655 : OAI22_X1 port map( A1 => n10842, A2 => n283, B1 => n5061, B2 => 
                           n131, ZN => n9570);
   U10656 : AOI22_X1 port map( A1 => n9491, A2 => n5062, B1 => n9492, B2 => 
                           n5063, ZN => n9568);
   U10657 : AOI22_X1 port map( A1 => n9493, A2 => n5064, B1 => n9494, B2 => 
                           n5065, ZN => n9567);
   U10658 : NAND3_X1 port map( A1 => n9571, A2 => n9572, A3 => n9573, ZN => 
                           n12204);
   U10659 : AOI221_X1 port map( B1 => n9488, B2 => n5069, C1 => n176, C2 => 
                           MEM_IN(20), A => n9574, ZN => n9573);
   U10660 : OAI22_X1 port map( A1 => n10841, A2 => n283, B1 => n5071, B2 => 
                           n131, ZN => n9574);
   U10661 : AOI22_X1 port map( A1 => n9491, A2 => n5072, B1 => n9492, B2 => 
                           n5073, ZN => n9572);
   U10662 : AOI22_X1 port map( A1 => n9493, A2 => n5074, B1 => n9494, B2 => 
                           n5075, ZN => n9571);
   U10663 : NAND3_X1 port map( A1 => n9575, A2 => n9576, A3 => n9577, ZN => 
                           n12203);
   U10664 : AOI221_X1 port map( B1 => n9488, B2 => n5079, C1 => n176, C2 => 
                           MEM_IN(21), A => n9578, ZN => n9577);
   U10665 : OAI22_X1 port map( A1 => n10840, A2 => n283, B1 => n5081, B2 => 
                           n131, ZN => n9578);
   U10666 : AOI22_X1 port map( A1 => n9491, A2 => n5082, B1 => n9492, B2 => 
                           n5083, ZN => n9576);
   U10667 : AOI22_X1 port map( A1 => n9493, A2 => n5084, B1 => n9494, B2 => 
                           n5085, ZN => n9575);
   U10668 : NAND3_X1 port map( A1 => n9579, A2 => n9580, A3 => n9581, ZN => 
                           n12202);
   U10669 : AOI221_X1 port map( B1 => n9488, B2 => n5089, C1 => n176, C2 => 
                           MEM_IN(22), A => n9582, ZN => n9581);
   U10670 : OAI22_X1 port map( A1 => n10839, A2 => n283, B1 => n5091, B2 => 
                           n131, ZN => n9582);
   U10671 : AOI22_X1 port map( A1 => n9491, A2 => n5092, B1 => n9492, B2 => 
                           n5093, ZN => n9580);
   U10672 : AOI22_X1 port map( A1 => n9493, A2 => n5094, B1 => n9494, B2 => 
                           n5095, ZN => n9579);
   U10673 : NAND3_X1 port map( A1 => n9583, A2 => n9584, A3 => n9585, ZN => 
                           n12201);
   U10674 : AOI221_X1 port map( B1 => n9488, B2 => n5099, C1 => n176, C2 => 
                           MEM_IN(23), A => n9586, ZN => n9585);
   U10675 : OAI22_X1 port map( A1 => n10838, A2 => n283, B1 => n5101, B2 => 
                           n131, ZN => n9586);
   U10676 : AOI22_X1 port map( A1 => n9491, A2 => n5102, B1 => n9492, B2 => 
                           n5103, ZN => n9584);
   U10677 : AOI22_X1 port map( A1 => n9493, A2 => n5104, B1 => n9494, B2 => 
                           n5105, ZN => n9583);
   U10678 : NAND3_X1 port map( A1 => n9587, A2 => n9588, A3 => n9589, ZN => 
                           n12200);
   U10679 : AOI221_X1 port map( B1 => n9488, B2 => n5109, C1 => n176, C2 => 
                           MEM_IN(24), A => n9590, ZN => n9589);
   U10680 : OAI22_X1 port map( A1 => n10837, A2 => n283, B1 => n5111, B2 => 
                           n131, ZN => n9590);
   U10681 : AOI22_X1 port map( A1 => n9491, A2 => n5112, B1 => n9492, B2 => 
                           n5113, ZN => n9588);
   U10682 : AOI22_X1 port map( A1 => n9493, A2 => n5114, B1 => n9494, B2 => 
                           n5115, ZN => n9587);
   U10683 : NAND3_X1 port map( A1 => n9591, A2 => n9592, A3 => n9593, ZN => 
                           n12199);
   U10684 : AOI221_X1 port map( B1 => n9488, B2 => n5119, C1 => n176, C2 => 
                           MEM_IN(25), A => n9594, ZN => n9593);
   U10685 : OAI22_X1 port map( A1 => n10836, A2 => n283, B1 => n5121, B2 => 
                           n131, ZN => n9594);
   U10686 : AOI22_X1 port map( A1 => n9491, A2 => n5122, B1 => n9492, B2 => 
                           n5123, ZN => n9592);
   U10687 : AOI22_X1 port map( A1 => n9493, A2 => n5124, B1 => n9494, B2 => 
                           n5125, ZN => n9591);
   U10688 : NAND3_X1 port map( A1 => n9595, A2 => n9596, A3 => n9597, ZN => 
                           n12198);
   U10689 : AOI221_X1 port map( B1 => n9488, B2 => n5129, C1 => n176, C2 => 
                           MEM_IN(26), A => n9598, ZN => n9597);
   U10690 : OAI22_X1 port map( A1 => n10835, A2 => n283, B1 => n5131, B2 => 
                           n131, ZN => n9598);
   U10691 : AOI22_X1 port map( A1 => n9491, A2 => n5132, B1 => n9492, B2 => 
                           n5133, ZN => n9596);
   U10692 : AOI22_X1 port map( A1 => n9493, A2 => n5134, B1 => n9494, B2 => 
                           n5135, ZN => n9595);
   U10693 : NAND3_X1 port map( A1 => n9599, A2 => n9600, A3 => n9601, ZN => 
                           n12197);
   U10694 : AOI221_X1 port map( B1 => n9488, B2 => n5139, C1 => n176, C2 => 
                           MEM_IN(27), A => n9602, ZN => n9601);
   U10695 : OAI22_X1 port map( A1 => n10834, A2 => n283, B1 => n5141, B2 => 
                           n131, ZN => n9602);
   U10696 : AOI22_X1 port map( A1 => n9491, A2 => n5142, B1 => n9492, B2 => 
                           n5143, ZN => n9600);
   U10697 : AOI22_X1 port map( A1 => n9493, A2 => n5144, B1 => n9494, B2 => 
                           n5145, ZN => n9599);
   U10698 : NAND3_X1 port map( A1 => n9603, A2 => n9604, A3 => n9605, ZN => 
                           n12196);
   U10699 : AOI221_X1 port map( B1 => n9488, B2 => n5149, C1 => n176, C2 => 
                           MEM_IN(28), A => n9606, ZN => n9605);
   U10700 : OAI22_X1 port map( A1 => n10833, A2 => n283, B1 => n5151, B2 => 
                           n131, ZN => n9606);
   U10701 : AOI22_X1 port map( A1 => n9491, A2 => n5152, B1 => n9492, B2 => 
                           n5153, ZN => n9604);
   U10702 : AOI22_X1 port map( A1 => n9493, A2 => n5154, B1 => n9494, B2 => 
                           n5155, ZN => n9603);
   U10703 : NAND3_X1 port map( A1 => n9607, A2 => n9608, A3 => n9609, ZN => 
                           n12195);
   U10704 : AOI221_X1 port map( B1 => n9488, B2 => n5159, C1 => n176, C2 => 
                           MEM_IN(29), A => n9610, ZN => n9609);
   U10705 : OAI22_X1 port map( A1 => n10832, A2 => n283, B1 => n5161, B2 => 
                           n131, ZN => n9610);
   U10706 : AOI22_X1 port map( A1 => n9491, A2 => n5162, B1 => n9492, B2 => 
                           n5163, ZN => n9608);
   U10707 : AOI22_X1 port map( A1 => n9493, A2 => n5164, B1 => n9494, B2 => 
                           n5165, ZN => n9607);
   U10708 : NAND3_X1 port map( A1 => n9611, A2 => n9612, A3 => n9613, ZN => 
                           n12194);
   U10709 : AOI221_X1 port map( B1 => n9488, B2 => n5169, C1 => n176, C2 => 
                           MEM_IN(30), A => n9614, ZN => n9613);
   U10710 : OAI22_X1 port map( A1 => n10831, A2 => n283, B1 => n5171, B2 => 
                           n131, ZN => n9614);
   U10711 : AOI22_X1 port map( A1 => n9491, A2 => n5172, B1 => n9492, B2 => 
                           n5173, ZN => n9612);
   U10712 : AOI22_X1 port map( A1 => n9493, A2 => n5174, B1 => n9494, B2 => 
                           n5175, ZN => n9611);
   U10713 : NAND3_X1 port map( A1 => n9615, A2 => n9616, A3 => n9617, ZN => 
                           n12193);
   U10714 : AOI221_X1 port map( B1 => n9488, B2 => n5179, C1 => n176, C2 => 
                           MEM_IN(31), A => n9618, ZN => n9617);
   U10715 : OAI22_X1 port map( A1 => n10830, A2 => n283, B1 => n5181, B2 => 
                           n131, ZN => n9618);
   U10716 : INV_X1 port map( A => n9622, ZN => n9621);
   U10717 : NAND2_X1 port map( A1 => n5206, A2 => n9476, ZN => n9474);
   U10718 : NAND3_X1 port map( A1 => n5206, A2 => n8745, A3 => n9189, ZN => 
                           n9476);
   U10719 : AOI22_X1 port map( A1 => n9491, A2 => n5191, B1 => n9492, B2 => 
                           n5192, ZN => n9616);
   U10720 : AOI22_X1 port map( A1 => n9493, A2 => n5195, B1 => n9494, B2 => 
                           n5196, ZN => n9615);
   U10721 : OAI22_X1 port map( A1 => n9622, A2 => n9620, B1 => n208, B2 => n282
                           , ZN => n9624);
   U10722 : NAND3_X1 port map( A1 => n208, A2 => n283, A3 => n8595, ZN => n9620
                           );
   U10723 : INV_X1 port map( A => n9619, ZN => n8595);
   U10724 : OAI22_X1 port map( A1 => n4786, A2 => n9626, B1 => n9627, B2 => 
                           n5204, ZN => n9490);
   U10725 : NOR2_X1 port map( A1 => n9619, A2 => n9622, ZN => n9627);
   U10726 : NAND3_X1 port map( A1 => n9336, A2 => n8745, A3 => n9628, ZN => 
                           n9619);
   U10727 : NOR3_X1 port map( A1 => n9629, A2 => RESET, A3 => n9186, ZN => 
                           n9626);
   U10728 : OAI22_X1 port map( A1 => n6076, A2 => n9043, B1 => n9336, B2 => 
                           n4787, ZN => n9629);
   U10729 : NAND2_X1 port map( A1 => n9630, A2 => n9631, ZN => n9622);
   U10730 : NOR2_X1 port map( A1 => n8745, A2 => n4787, ZN => n9186);
   U10731 : NAND2_X1 port map( A1 => n8895, A2 => n6079, ZN => n8745);
   U10732 : NAND3_X1 port map( A1 => n9632, A2 => n9633, A3 => n9634, ZN => 
                           n12192);
   U10733 : AOI221_X1 port map( B1 => n9635, B2 => n4863, C1 => n177, C2 => 
                           MEM_IN(0), A => n9636, ZN => n9634);
   U10734 : OAI22_X1 port map( A1 => n10829, A2 => n269, B1 => n4867, B2 => 
                           n128, ZN => n9636);
   U10735 : AOI22_X1 port map( A1 => n9638, A2 => n4869, B1 => n9639, B2 => 
                           n4871, ZN => n9633);
   U10736 : AOI22_X1 port map( A1 => n9640, A2 => n4873, B1 => n9641, B2 => 
                           n4875, ZN => n9632);
   U10737 : NAND3_X1 port map( A1 => n9642, A2 => n9643, A3 => n9644, ZN => 
                           n12191);
   U10738 : AOI221_X1 port map( B1 => n9635, B2 => n4879, C1 => n177, C2 => 
                           MEM_IN(1), A => n9645, ZN => n9644);
   U10739 : OAI22_X1 port map( A1 => n10828, A2 => n269, B1 => n4881, B2 => 
                           n128, ZN => n9645);
   U10740 : AOI22_X1 port map( A1 => n9638, A2 => n4882, B1 => n9639, B2 => 
                           n4883, ZN => n9643);
   U10741 : AOI22_X1 port map( A1 => n9640, A2 => n4884, B1 => n9641, B2 => 
                           n4885, ZN => n9642);
   U10742 : NAND3_X1 port map( A1 => n9646, A2 => n9647, A3 => n9648, ZN => 
                           n12190);
   U10743 : AOI221_X1 port map( B1 => n9635, B2 => n4889, C1 => n177, C2 => 
                           MEM_IN(2), A => n9649, ZN => n9648);
   U10744 : OAI22_X1 port map( A1 => n10827, A2 => n269, B1 => n4891, B2 => 
                           n128, ZN => n9649);
   U10745 : AOI22_X1 port map( A1 => n9638, A2 => n4892, B1 => n9639, B2 => 
                           n4893, ZN => n9647);
   U10746 : AOI22_X1 port map( A1 => n9640, A2 => n4894, B1 => n9641, B2 => 
                           n4895, ZN => n9646);
   U10747 : NAND3_X1 port map( A1 => n9650, A2 => n9651, A3 => n9652, ZN => 
                           n12189);
   U10748 : AOI221_X1 port map( B1 => n9635, B2 => n4899, C1 => n177, C2 => 
                           MEM_IN(3), A => n9653, ZN => n9652);
   U10749 : OAI22_X1 port map( A1 => n10826, A2 => n269, B1 => n4901, B2 => 
                           n128, ZN => n9653);
   U10750 : AOI22_X1 port map( A1 => n9638, A2 => n4902, B1 => n9639, B2 => 
                           n4903, ZN => n9651);
   U10751 : AOI22_X1 port map( A1 => n9640, A2 => n4904, B1 => n9641, B2 => 
                           n4905, ZN => n9650);
   U10752 : NAND3_X1 port map( A1 => n9654, A2 => n9655, A3 => n9656, ZN => 
                           n12188);
   U10753 : AOI221_X1 port map( B1 => n9635, B2 => n4909, C1 => n177, C2 => 
                           MEM_IN(4), A => n9657, ZN => n9656);
   U10754 : OAI22_X1 port map( A1 => n10825, A2 => n269, B1 => n4911, B2 => 
                           n128, ZN => n9657);
   U10755 : AOI22_X1 port map( A1 => n9638, A2 => n4912, B1 => n9639, B2 => 
                           n4913, ZN => n9655);
   U10756 : AOI22_X1 port map( A1 => n9640, A2 => n4914, B1 => n9641, B2 => 
                           n4915, ZN => n9654);
   U10757 : NAND3_X1 port map( A1 => n9658, A2 => n9659, A3 => n9660, ZN => 
                           n12187);
   U10758 : AOI221_X1 port map( B1 => n9635, B2 => n4919, C1 => n177, C2 => 
                           MEM_IN(5), A => n9661, ZN => n9660);
   U10759 : OAI22_X1 port map( A1 => n10824, A2 => n269, B1 => n4921, B2 => 
                           n128, ZN => n9661);
   U10760 : AOI22_X1 port map( A1 => n9638, A2 => n4922, B1 => n9639, B2 => 
                           n4923, ZN => n9659);
   U10761 : AOI22_X1 port map( A1 => n9640, A2 => n4924, B1 => n9641, B2 => 
                           n4925, ZN => n9658);
   U10762 : NAND3_X1 port map( A1 => n9662, A2 => n9663, A3 => n9664, ZN => 
                           n12186);
   U10763 : AOI221_X1 port map( B1 => n9635, B2 => n4929, C1 => n177, C2 => 
                           MEM_IN(6), A => n9665, ZN => n9664);
   U10764 : OAI22_X1 port map( A1 => n10823, A2 => n269, B1 => n4931, B2 => 
                           n128, ZN => n9665);
   U10765 : AOI22_X1 port map( A1 => n9638, A2 => n4932, B1 => n9639, B2 => 
                           n4933, ZN => n9663);
   U10766 : AOI22_X1 port map( A1 => n9640, A2 => n4934, B1 => n9641, B2 => 
                           n4935, ZN => n9662);
   U10767 : NAND3_X1 port map( A1 => n9666, A2 => n9667, A3 => n9668, ZN => 
                           n12185);
   U10768 : AOI221_X1 port map( B1 => n9635, B2 => n4939, C1 => n177, C2 => 
                           MEM_IN(7), A => n9669, ZN => n9668);
   U10769 : OAI22_X1 port map( A1 => n10822, A2 => n269, B1 => n4941, B2 => 
                           n128, ZN => n9669);
   U10770 : AOI22_X1 port map( A1 => n9638, A2 => n4942, B1 => n9639, B2 => 
                           n4943, ZN => n9667);
   U10771 : AOI22_X1 port map( A1 => n9640, A2 => n4944, B1 => n9641, B2 => 
                           n4945, ZN => n9666);
   U10772 : NAND3_X1 port map( A1 => n9670, A2 => n9671, A3 => n9672, ZN => 
                           n12184);
   U10773 : AOI221_X1 port map( B1 => n9635, B2 => n4949, C1 => n177, C2 => 
                           MEM_IN(8), A => n9673, ZN => n9672);
   U10774 : OAI22_X1 port map( A1 => n10821, A2 => n269, B1 => n4951, B2 => 
                           n128, ZN => n9673);
   U10775 : AOI22_X1 port map( A1 => n9638, A2 => n4952, B1 => n9639, B2 => 
                           n4953, ZN => n9671);
   U10776 : AOI22_X1 port map( A1 => n9640, A2 => n4954, B1 => n9641, B2 => 
                           n4955, ZN => n9670);
   U10777 : NAND3_X1 port map( A1 => n9674, A2 => n9675, A3 => n9676, ZN => 
                           n12183);
   U10778 : AOI221_X1 port map( B1 => n9635, B2 => n4959, C1 => n177, C2 => 
                           MEM_IN(9), A => n9677, ZN => n9676);
   U10779 : OAI22_X1 port map( A1 => n10820, A2 => n269, B1 => n4961, B2 => 
                           n128, ZN => n9677);
   U10780 : AOI22_X1 port map( A1 => n9638, A2 => n4962, B1 => n9639, B2 => 
                           n4963, ZN => n9675);
   U10781 : AOI22_X1 port map( A1 => n9640, A2 => n4964, B1 => n9641, B2 => 
                           n4965, ZN => n9674);
   U10782 : NAND3_X1 port map( A1 => n9678, A2 => n9679, A3 => n9680, ZN => 
                           n12182);
   U10783 : AOI221_X1 port map( B1 => n9635, B2 => n4969, C1 => n177, C2 => 
                           MEM_IN(10), A => n9681, ZN => n9680);
   U10784 : OAI22_X1 port map( A1 => n10819, A2 => n269, B1 => n4971, B2 => 
                           n128, ZN => n9681);
   U10785 : AOI22_X1 port map( A1 => n9638, A2 => n4972, B1 => n9639, B2 => 
                           n4973, ZN => n9679);
   U10786 : AOI22_X1 port map( A1 => n9640, A2 => n4974, B1 => n9641, B2 => 
                           n4975, ZN => n9678);
   U10787 : NAND3_X1 port map( A1 => n9682, A2 => n9683, A3 => n9684, ZN => 
                           n12181);
   U10788 : AOI221_X1 port map( B1 => n9635, B2 => n4979, C1 => n177, C2 => 
                           MEM_IN(11), A => n9685, ZN => n9684);
   U10789 : OAI22_X1 port map( A1 => n10818, A2 => n269, B1 => n4981, B2 => 
                           n128, ZN => n9685);
   U10790 : AOI22_X1 port map( A1 => n9638, A2 => n4982, B1 => n9639, B2 => 
                           n4983, ZN => n9683);
   U10791 : AOI22_X1 port map( A1 => n9640, A2 => n4984, B1 => n9641, B2 => 
                           n4985, ZN => n9682);
   U10792 : NAND3_X1 port map( A1 => n9686, A2 => n9687, A3 => n9688, ZN => 
                           n12180);
   U10793 : AOI221_X1 port map( B1 => n9635, B2 => n4989, C1 => n177, C2 => 
                           MEM_IN(12), A => n9689, ZN => n9688);
   U10794 : OAI22_X1 port map( A1 => n10817, A2 => n269, B1 => n4991, B2 => 
                           n128, ZN => n9689);
   U10795 : AOI22_X1 port map( A1 => n9638, A2 => n4992, B1 => n9639, B2 => 
                           n4993, ZN => n9687);
   U10796 : AOI22_X1 port map( A1 => n9640, A2 => n4994, B1 => n9641, B2 => 
                           n4995, ZN => n9686);
   U10797 : NAND3_X1 port map( A1 => n9690, A2 => n9691, A3 => n9692, ZN => 
                           n12179);
   U10798 : AOI221_X1 port map( B1 => n9635, B2 => n4999, C1 => n177, C2 => 
                           MEM_IN(13), A => n9693, ZN => n9692);
   U10799 : OAI22_X1 port map( A1 => n10816, A2 => n269, B1 => n5001, B2 => 
                           n128, ZN => n9693);
   U10800 : AOI22_X1 port map( A1 => n9638, A2 => n5002, B1 => n9639, B2 => 
                           n5003, ZN => n9691);
   U10801 : AOI22_X1 port map( A1 => n9640, A2 => n5004, B1 => n9641, B2 => 
                           n5005, ZN => n9690);
   U10802 : NAND3_X1 port map( A1 => n9694, A2 => n9695, A3 => n9696, ZN => 
                           n12178);
   U10803 : AOI221_X1 port map( B1 => n9635, B2 => n5009, C1 => n177, C2 => 
                           MEM_IN(14), A => n9697, ZN => n9696);
   U10804 : OAI22_X1 port map( A1 => n10815, A2 => n269, B1 => n5011, B2 => 
                           n128, ZN => n9697);
   U10805 : AOI22_X1 port map( A1 => n9638, A2 => n5012, B1 => n9639, B2 => 
                           n5013, ZN => n9695);
   U10806 : AOI22_X1 port map( A1 => n9640, A2 => n5014, B1 => n9641, B2 => 
                           n5015, ZN => n9694);
   U10807 : NAND3_X1 port map( A1 => n9698, A2 => n9699, A3 => n9700, ZN => 
                           n12177);
   U10808 : AOI221_X1 port map( B1 => n9635, B2 => n5019, C1 => n177, C2 => 
                           MEM_IN(15), A => n9701, ZN => n9700);
   U10809 : OAI22_X1 port map( A1 => n10814, A2 => n269, B1 => n5021, B2 => 
                           n128, ZN => n9701);
   U10810 : AOI22_X1 port map( A1 => n9638, A2 => n5022, B1 => n9639, B2 => 
                           n5023, ZN => n9699);
   U10811 : AOI22_X1 port map( A1 => n9640, A2 => n5024, B1 => n9641, B2 => 
                           n5025, ZN => n9698);
   U10812 : NAND3_X1 port map( A1 => n9702, A2 => n9703, A3 => n9704, ZN => 
                           n12176);
   U10813 : AOI221_X1 port map( B1 => n9635, B2 => n5029, C1 => n177, C2 => 
                           MEM_IN(16), A => n9705, ZN => n9704);
   U10814 : OAI22_X1 port map( A1 => n10813, A2 => n269, B1 => n5031, B2 => 
                           n128, ZN => n9705);
   U10815 : AOI22_X1 port map( A1 => n9638, A2 => n5032, B1 => n9639, B2 => 
                           n5033, ZN => n9703);
   U10816 : AOI22_X1 port map( A1 => n9640, A2 => n5034, B1 => n9641, B2 => 
                           n5035, ZN => n9702);
   U10817 : NAND3_X1 port map( A1 => n9706, A2 => n9707, A3 => n9708, ZN => 
                           n12175);
   U10818 : AOI221_X1 port map( B1 => n9635, B2 => n5039, C1 => n177, C2 => 
                           MEM_IN(17), A => n9709, ZN => n9708);
   U10819 : OAI22_X1 port map( A1 => n10812, A2 => n269, B1 => n5041, B2 => 
                           n128, ZN => n9709);
   U10820 : AOI22_X1 port map( A1 => n9638, A2 => n5042, B1 => n9639, B2 => 
                           n5043, ZN => n9707);
   U10821 : AOI22_X1 port map( A1 => n9640, A2 => n5044, B1 => n9641, B2 => 
                           n5045, ZN => n9706);
   U10822 : NAND3_X1 port map( A1 => n9710, A2 => n9711, A3 => n9712, ZN => 
                           n12174);
   U10823 : AOI221_X1 port map( B1 => n9635, B2 => n5049, C1 => n177, C2 => 
                           MEM_IN(18), A => n9713, ZN => n9712);
   U10824 : OAI22_X1 port map( A1 => n10811, A2 => n269, B1 => n5051, B2 => 
                           n128, ZN => n9713);
   U10825 : AOI22_X1 port map( A1 => n9638, A2 => n5052, B1 => n9639, B2 => 
                           n5053, ZN => n9711);
   U10826 : AOI22_X1 port map( A1 => n9640, A2 => n5054, B1 => n9641, B2 => 
                           n5055, ZN => n9710);
   U10827 : NAND3_X1 port map( A1 => n9714, A2 => n9715, A3 => n9716, ZN => 
                           n12173);
   U10828 : AOI221_X1 port map( B1 => n9635, B2 => n5059, C1 => n177, C2 => 
                           MEM_IN(19), A => n9717, ZN => n9716);
   U10829 : OAI22_X1 port map( A1 => n10810, A2 => n269, B1 => n5061, B2 => 
                           n128, ZN => n9717);
   U10830 : AOI22_X1 port map( A1 => n9638, A2 => n5062, B1 => n9639, B2 => 
                           n5063, ZN => n9715);
   U10831 : AOI22_X1 port map( A1 => n9640, A2 => n5064, B1 => n9641, B2 => 
                           n5065, ZN => n9714);
   U10832 : NAND3_X1 port map( A1 => n9718, A2 => n9719, A3 => n9720, ZN => 
                           n12172);
   U10833 : AOI221_X1 port map( B1 => n9635, B2 => n5069, C1 => n177, C2 => 
                           MEM_IN(20), A => n9721, ZN => n9720);
   U10834 : OAI22_X1 port map( A1 => n10809, A2 => n269, B1 => n5071, B2 => 
                           n128, ZN => n9721);
   U10835 : AOI22_X1 port map( A1 => n9638, A2 => n5072, B1 => n9639, B2 => 
                           n5073, ZN => n9719);
   U10836 : AOI22_X1 port map( A1 => n9640, A2 => n5074, B1 => n9641, B2 => 
                           n5075, ZN => n9718);
   U10837 : NAND3_X1 port map( A1 => n9722, A2 => n9723, A3 => n9724, ZN => 
                           n12171);
   U10838 : AOI221_X1 port map( B1 => n9635, B2 => n5079, C1 => n177, C2 => 
                           MEM_IN(21), A => n9725, ZN => n9724);
   U10839 : OAI22_X1 port map( A1 => n10808, A2 => n269, B1 => n5081, B2 => 
                           n128, ZN => n9725);
   U10840 : AOI22_X1 port map( A1 => n9638, A2 => n5082, B1 => n9639, B2 => 
                           n5083, ZN => n9723);
   U10841 : AOI22_X1 port map( A1 => n9640, A2 => n5084, B1 => n9641, B2 => 
                           n5085, ZN => n9722);
   U10842 : NAND3_X1 port map( A1 => n9726, A2 => n9727, A3 => n9728, ZN => 
                           n12170);
   U10843 : AOI221_X1 port map( B1 => n9635, B2 => n5089, C1 => n177, C2 => 
                           MEM_IN(22), A => n9729, ZN => n9728);
   U10844 : OAI22_X1 port map( A1 => n10807, A2 => n269, B1 => n5091, B2 => 
                           n128, ZN => n9729);
   U10845 : AOI22_X1 port map( A1 => n9638, A2 => n5092, B1 => n9639, B2 => 
                           n5093, ZN => n9727);
   U10846 : AOI22_X1 port map( A1 => n9640, A2 => n5094, B1 => n9641, B2 => 
                           n5095, ZN => n9726);
   U10847 : NAND3_X1 port map( A1 => n9730, A2 => n9731, A3 => n9732, ZN => 
                           n12169);
   U10848 : AOI221_X1 port map( B1 => n9635, B2 => n5099, C1 => n177, C2 => 
                           MEM_IN(23), A => n9733, ZN => n9732);
   U10849 : OAI22_X1 port map( A1 => n10806, A2 => n269, B1 => n5101, B2 => 
                           n128, ZN => n9733);
   U10850 : AOI22_X1 port map( A1 => n9638, A2 => n5102, B1 => n9639, B2 => 
                           n5103, ZN => n9731);
   U10851 : AOI22_X1 port map( A1 => n9640, A2 => n5104, B1 => n9641, B2 => 
                           n5105, ZN => n9730);
   U10852 : NAND3_X1 port map( A1 => n9734, A2 => n9735, A3 => n9736, ZN => 
                           n12168);
   U10853 : AOI221_X1 port map( B1 => n9635, B2 => n5109, C1 => n177, C2 => 
                           MEM_IN(24), A => n9737, ZN => n9736);
   U10854 : OAI22_X1 port map( A1 => n10805, A2 => n269, B1 => n5111, B2 => 
                           n128, ZN => n9737);
   U10855 : AOI22_X1 port map( A1 => n9638, A2 => n5112, B1 => n9639, B2 => 
                           n5113, ZN => n9735);
   U10856 : AOI22_X1 port map( A1 => n9640, A2 => n5114, B1 => n9641, B2 => 
                           n5115, ZN => n9734);
   U10857 : NAND3_X1 port map( A1 => n9738, A2 => n9739, A3 => n9740, ZN => 
                           n12167);
   U10858 : AOI221_X1 port map( B1 => n9635, B2 => n5119, C1 => n177, C2 => 
                           MEM_IN(25), A => n9741, ZN => n9740);
   U10859 : OAI22_X1 port map( A1 => n10804, A2 => n269, B1 => n5121, B2 => 
                           n128, ZN => n9741);
   U10860 : AOI22_X1 port map( A1 => n9638, A2 => n5122, B1 => n9639, B2 => 
                           n5123, ZN => n9739);
   U10861 : AOI22_X1 port map( A1 => n9640, A2 => n5124, B1 => n9641, B2 => 
                           n5125, ZN => n9738);
   U10862 : NAND3_X1 port map( A1 => n9742, A2 => n9743, A3 => n9744, ZN => 
                           n12166);
   U10863 : AOI221_X1 port map( B1 => n9635, B2 => n5129, C1 => n177, C2 => 
                           MEM_IN(26), A => n9745, ZN => n9744);
   U10864 : OAI22_X1 port map( A1 => n10803, A2 => n269, B1 => n5131, B2 => 
                           n128, ZN => n9745);
   U10865 : AOI22_X1 port map( A1 => n9638, A2 => n5132, B1 => n9639, B2 => 
                           n5133, ZN => n9743);
   U10866 : AOI22_X1 port map( A1 => n9640, A2 => n5134, B1 => n9641, B2 => 
                           n5135, ZN => n9742);
   U10867 : NAND3_X1 port map( A1 => n9746, A2 => n9747, A3 => n9748, ZN => 
                           n12165);
   U10868 : AOI221_X1 port map( B1 => n9635, B2 => n5139, C1 => n177, C2 => 
                           MEM_IN(27), A => n9749, ZN => n9748);
   U10869 : OAI22_X1 port map( A1 => n10802, A2 => n269, B1 => n5141, B2 => 
                           n128, ZN => n9749);
   U10870 : AOI22_X1 port map( A1 => n9638, A2 => n5142, B1 => n9639, B2 => 
                           n5143, ZN => n9747);
   U10871 : AOI22_X1 port map( A1 => n9640, A2 => n5144, B1 => n9641, B2 => 
                           n5145, ZN => n9746);
   U10872 : NAND3_X1 port map( A1 => n9750, A2 => n9751, A3 => n9752, ZN => 
                           n12164);
   U10873 : AOI221_X1 port map( B1 => n9635, B2 => n5149, C1 => n177, C2 => 
                           MEM_IN(28), A => n9753, ZN => n9752);
   U10874 : OAI22_X1 port map( A1 => n10801, A2 => n269, B1 => n5151, B2 => 
                           n128, ZN => n9753);
   U10875 : AOI22_X1 port map( A1 => n9638, A2 => n5152, B1 => n9639, B2 => 
                           n5153, ZN => n9751);
   U10876 : AOI22_X1 port map( A1 => n9640, A2 => n5154, B1 => n9641, B2 => 
                           n5155, ZN => n9750);
   U10877 : NAND3_X1 port map( A1 => n9754, A2 => n9755, A3 => n9756, ZN => 
                           n12163);
   U10878 : AOI221_X1 port map( B1 => n9635, B2 => n5159, C1 => n177, C2 => 
                           MEM_IN(29), A => n9757, ZN => n9756);
   U10879 : OAI22_X1 port map( A1 => n10800, A2 => n269, B1 => n5161, B2 => 
                           n128, ZN => n9757);
   U10880 : AOI22_X1 port map( A1 => n9638, A2 => n5162, B1 => n9639, B2 => 
                           n5163, ZN => n9755);
   U10881 : AOI22_X1 port map( A1 => n9640, A2 => n5164, B1 => n9641, B2 => 
                           n5165, ZN => n9754);
   U10882 : NAND3_X1 port map( A1 => n9758, A2 => n9759, A3 => n9760, ZN => 
                           n12162);
   U10883 : AOI221_X1 port map( B1 => n9635, B2 => n5169, C1 => n177, C2 => 
                           MEM_IN(30), A => n9761, ZN => n9760);
   U10884 : OAI22_X1 port map( A1 => n10799, A2 => n269, B1 => n5171, B2 => 
                           n128, ZN => n9761);
   U10885 : AOI22_X1 port map( A1 => n9638, A2 => n5172, B1 => n9639, B2 => 
                           n5173, ZN => n9759);
   U10886 : AOI22_X1 port map( A1 => n9640, A2 => n5174, B1 => n9641, B2 => 
                           n5175, ZN => n9758);
   U10887 : NAND3_X1 port map( A1 => n9762, A2 => n9763, A3 => n9764, ZN => 
                           n12161);
   U10888 : AOI221_X1 port map( B1 => n9635, B2 => n5179, C1 => n177, C2 => 
                           MEM_IN(31), A => n9765, ZN => n9764);
   U10889 : OAI22_X1 port map( A1 => n10798, A2 => n269, B1 => n5181, B2 => 
                           n128, ZN => n9765);
   U10890 : INV_X1 port map( A => n9769, ZN => n9768);
   U10891 : AOI22_X1 port map( A1 => n9638, A2 => n5191, B1 => n9639, B2 => 
                           n5192, ZN => n9763);
   U10892 : AOI22_X1 port map( A1 => n9640, A2 => n5195, B1 => n9641, B2 => 
                           n5196, ZN => n9762);
   U10893 : OAI22_X1 port map( A1 => n9769, A2 => n9767, B1 => n208, B2 => n268
                           , ZN => n9771);
   U10894 : NAND3_X1 port map( A1 => n208, A2 => n269, A3 => n8744, ZN => n9767
                           );
   U10895 : INV_X1 port map( A => n9766, ZN => n8744);
   U10896 : OAI22_X1 port map( A1 => n4786, A2 => n9773, B1 => n9774, B2 => 
                           n5204, ZN => n9637);
   U10897 : NOR2_X1 port map( A1 => n9766, A2 => n9769, ZN => n9774);
   U10898 : NAND2_X1 port map( A1 => n9775, A2 => n9336, ZN => n9766);
   U10899 : INV_X1 port map( A => n9776, ZN => n9336);
   U10900 : INV_X1 port map( A => n9777, ZN => n9773);
   U10901 : OAI211_X1 port map( C1 => n9043, C2 => n8594, A => n9770, B => 
                           n5368, ZN => n9777);
   U10902 : AOI21_X1 port map( B1 => n9776, B2 => n5206, A => n9772, ZN => 
                           n9770);
   U10903 : NAND2_X1 port map( A1 => n9189, A2 => n9192, ZN => n9776);
   U10904 : AND2_X1 port map( A1 => n9045, A2 => n8894, ZN => n9189);
   U10905 : NAND2_X1 port map( A1 => n9778, A2 => n9779, ZN => n9769);
   U10906 : NOR2_X1 port map( A1 => n8894, A2 => n4787, ZN => n9333);
   U10907 : NAND2_X1 port map( A1 => n8895, A2 => n6228, ZN => n8894);
   U10908 : NAND3_X1 port map( A1 => n9780, A2 => n9781, A3 => n9782, ZN => 
                           n12160);
   U10909 : AOI221_X1 port map( B1 => n9783, B2 => n4863, C1 => n174, C2 => 
                           MEM_IN(0), A => n9784, ZN => n9782);
   U10910 : OAI22_X1 port map( A1 => n10797, A2 => n257, B1 => n4867, B2 => 
                           n129, ZN => n9784);
   U10911 : AOI22_X1 port map( A1 => n9786, A2 => n4869, B1 => n9787, B2 => 
                           n4871, ZN => n9781);
   U10912 : AOI22_X1 port map( A1 => n238, A2 => n4873, B1 => n9788, B2 => 
                           n4875, ZN => n9780);
   U10913 : NAND3_X1 port map( A1 => n9789, A2 => n9790, A3 => n9791, ZN => 
                           n12159);
   U10914 : AOI221_X1 port map( B1 => n9783, B2 => n4879, C1 => n174, C2 => 
                           MEM_IN(1), A => n9792, ZN => n9791);
   U10915 : OAI22_X1 port map( A1 => n10796, A2 => n257, B1 => n4881, B2 => 
                           n129, ZN => n9792);
   U10916 : AOI22_X1 port map( A1 => n9786, A2 => n4882, B1 => n9787, B2 => 
                           n4883, ZN => n9790);
   U10917 : AOI22_X1 port map( A1 => n238, A2 => n4884, B1 => n9788, B2 => 
                           n4885, ZN => n9789);
   U10918 : NAND3_X1 port map( A1 => n9793, A2 => n9794, A3 => n9795, ZN => 
                           n12158);
   U10919 : AOI221_X1 port map( B1 => n9783, B2 => n4889, C1 => n174, C2 => 
                           MEM_IN(2), A => n9796, ZN => n9795);
   U10920 : OAI22_X1 port map( A1 => n10795, A2 => n257, B1 => n4891, B2 => 
                           n129, ZN => n9796);
   U10921 : AOI22_X1 port map( A1 => n9786, A2 => n4892, B1 => n9787, B2 => 
                           n4893, ZN => n9794);
   U10922 : AOI22_X1 port map( A1 => n238, A2 => n4894, B1 => n9788, B2 => 
                           n4895, ZN => n9793);
   U10923 : NAND3_X1 port map( A1 => n9797, A2 => n9798, A3 => n9799, ZN => 
                           n12157);
   U10924 : AOI221_X1 port map( B1 => n9783, B2 => n4899, C1 => n174, C2 => 
                           MEM_IN(3), A => n9800, ZN => n9799);
   U10925 : OAI22_X1 port map( A1 => n10794, A2 => n257, B1 => n4901, B2 => 
                           n129, ZN => n9800);
   U10926 : AOI22_X1 port map( A1 => n9786, A2 => n4902, B1 => n9787, B2 => 
                           n4903, ZN => n9798);
   U10927 : AOI22_X1 port map( A1 => n238, A2 => n4904, B1 => n9788, B2 => 
                           n4905, ZN => n9797);
   U10928 : NAND3_X1 port map( A1 => n9801, A2 => n9802, A3 => n9803, ZN => 
                           n12156);
   U10929 : AOI221_X1 port map( B1 => n9783, B2 => n4909, C1 => n174, C2 => 
                           MEM_IN(4), A => n9804, ZN => n9803);
   U10930 : OAI22_X1 port map( A1 => n10793, A2 => n257, B1 => n4911, B2 => 
                           n129, ZN => n9804);
   U10931 : AOI22_X1 port map( A1 => n9786, A2 => n4912, B1 => n9787, B2 => 
                           n4913, ZN => n9802);
   U10932 : AOI22_X1 port map( A1 => n238, A2 => n4914, B1 => n9788, B2 => 
                           n4915, ZN => n9801);
   U10933 : NAND3_X1 port map( A1 => n9805, A2 => n9806, A3 => n9807, ZN => 
                           n12155);
   U10934 : AOI221_X1 port map( B1 => n9783, B2 => n4919, C1 => n174, C2 => 
                           MEM_IN(5), A => n9808, ZN => n9807);
   U10935 : OAI22_X1 port map( A1 => n10792, A2 => n257, B1 => n4921, B2 => 
                           n129, ZN => n9808);
   U10936 : AOI22_X1 port map( A1 => n9786, A2 => n4922, B1 => n9787, B2 => 
                           n4923, ZN => n9806);
   U10937 : AOI22_X1 port map( A1 => n238, A2 => n4924, B1 => n9788, B2 => 
                           n4925, ZN => n9805);
   U10938 : NAND3_X1 port map( A1 => n9809, A2 => n9810, A3 => n9811, ZN => 
                           n12154);
   U10939 : AOI221_X1 port map( B1 => n9783, B2 => n4929, C1 => n174, C2 => 
                           MEM_IN(6), A => n9812, ZN => n9811);
   U10940 : OAI22_X1 port map( A1 => n10791, A2 => n257, B1 => n4931, B2 => 
                           n129, ZN => n9812);
   U10941 : AOI22_X1 port map( A1 => n9786, A2 => n4932, B1 => n9787, B2 => 
                           n4933, ZN => n9810);
   U10942 : AOI22_X1 port map( A1 => n238, A2 => n4934, B1 => n9788, B2 => 
                           n4935, ZN => n9809);
   U10943 : NAND3_X1 port map( A1 => n9813, A2 => n9814, A3 => n9815, ZN => 
                           n12153);
   U10944 : AOI221_X1 port map( B1 => n9783, B2 => n4939, C1 => n174, C2 => 
                           MEM_IN(7), A => n9816, ZN => n9815);
   U10945 : OAI22_X1 port map( A1 => n10790, A2 => n257, B1 => n4941, B2 => 
                           n129, ZN => n9816);
   U10946 : AOI22_X1 port map( A1 => n9786, A2 => n4942, B1 => n9787, B2 => 
                           n4943, ZN => n9814);
   U10947 : AOI22_X1 port map( A1 => n238, A2 => n4944, B1 => n9788, B2 => 
                           n4945, ZN => n9813);
   U10948 : NAND3_X1 port map( A1 => n9817, A2 => n9818, A3 => n9819, ZN => 
                           n12152);
   U10949 : AOI221_X1 port map( B1 => n9783, B2 => n4949, C1 => n174, C2 => 
                           MEM_IN(8), A => n9820, ZN => n9819);
   U10950 : OAI22_X1 port map( A1 => n10789, A2 => n257, B1 => n4951, B2 => 
                           n129, ZN => n9820);
   U10951 : AOI22_X1 port map( A1 => n9786, A2 => n4952, B1 => n9787, B2 => 
                           n4953, ZN => n9818);
   U10952 : AOI22_X1 port map( A1 => n238, A2 => n4954, B1 => n9788, B2 => 
                           n4955, ZN => n9817);
   U10953 : NAND3_X1 port map( A1 => n9821, A2 => n9822, A3 => n9823, ZN => 
                           n12151);
   U10954 : AOI221_X1 port map( B1 => n9783, B2 => n4959, C1 => n174, C2 => 
                           MEM_IN(9), A => n9824, ZN => n9823);
   U10955 : OAI22_X1 port map( A1 => n10788, A2 => n257, B1 => n4961, B2 => 
                           n129, ZN => n9824);
   U10956 : AOI22_X1 port map( A1 => n9786, A2 => n4962, B1 => n9787, B2 => 
                           n4963, ZN => n9822);
   U10957 : AOI22_X1 port map( A1 => n238, A2 => n4964, B1 => n9788, B2 => 
                           n4965, ZN => n9821);
   U10958 : NAND3_X1 port map( A1 => n9825, A2 => n9826, A3 => n9827, ZN => 
                           n12150);
   U10959 : AOI221_X1 port map( B1 => n9783, B2 => n4969, C1 => n174, C2 => 
                           MEM_IN(10), A => n9828, ZN => n9827);
   U10960 : OAI22_X1 port map( A1 => n10787, A2 => n257, B1 => n4971, B2 => 
                           n129, ZN => n9828);
   U10961 : AOI22_X1 port map( A1 => n9786, A2 => n4972, B1 => n9787, B2 => 
                           n4973, ZN => n9826);
   U10962 : AOI22_X1 port map( A1 => n238, A2 => n4974, B1 => n9788, B2 => 
                           n4975, ZN => n9825);
   U10963 : NAND3_X1 port map( A1 => n9829, A2 => n9830, A3 => n9831, ZN => 
                           n12149);
   U10964 : AOI221_X1 port map( B1 => n9783, B2 => n4979, C1 => n174, C2 => 
                           MEM_IN(11), A => n9832, ZN => n9831);
   U10965 : OAI22_X1 port map( A1 => n10786, A2 => n257, B1 => n4981, B2 => 
                           n129, ZN => n9832);
   U10966 : AOI22_X1 port map( A1 => n9786, A2 => n4982, B1 => n9787, B2 => 
                           n4983, ZN => n9830);
   U10967 : AOI22_X1 port map( A1 => n238, A2 => n4984, B1 => n9788, B2 => 
                           n4985, ZN => n9829);
   U10968 : NAND3_X1 port map( A1 => n9833, A2 => n9834, A3 => n9835, ZN => 
                           n12148);
   U10969 : AOI221_X1 port map( B1 => n9783, B2 => n4989, C1 => n174, C2 => 
                           MEM_IN(12), A => n9836, ZN => n9835);
   U10970 : OAI22_X1 port map( A1 => n10785, A2 => n257, B1 => n4991, B2 => 
                           n129, ZN => n9836);
   U10971 : AOI22_X1 port map( A1 => n9786, A2 => n4992, B1 => n9787, B2 => 
                           n4993, ZN => n9834);
   U10972 : AOI22_X1 port map( A1 => n238, A2 => n4994, B1 => n9788, B2 => 
                           n4995, ZN => n9833);
   U10973 : NAND3_X1 port map( A1 => n9837, A2 => n9838, A3 => n9839, ZN => 
                           n12147);
   U10974 : AOI221_X1 port map( B1 => n9783, B2 => n4999, C1 => n174, C2 => 
                           MEM_IN(13), A => n9840, ZN => n9839);
   U10975 : OAI22_X1 port map( A1 => n10784, A2 => n257, B1 => n5001, B2 => 
                           n129, ZN => n9840);
   U10976 : AOI22_X1 port map( A1 => n9786, A2 => n5002, B1 => n9787, B2 => 
                           n5003, ZN => n9838);
   U10977 : AOI22_X1 port map( A1 => n238, A2 => n5004, B1 => n9788, B2 => 
                           n5005, ZN => n9837);
   U10978 : NAND3_X1 port map( A1 => n9841, A2 => n9842, A3 => n9843, ZN => 
                           n12146);
   U10979 : AOI221_X1 port map( B1 => n9783, B2 => n5009, C1 => n174, C2 => 
                           MEM_IN(14), A => n9844, ZN => n9843);
   U10980 : OAI22_X1 port map( A1 => n10783, A2 => n257, B1 => n5011, B2 => 
                           n129, ZN => n9844);
   U10981 : AOI22_X1 port map( A1 => n9786, A2 => n5012, B1 => n9787, B2 => 
                           n5013, ZN => n9842);
   U10982 : AOI22_X1 port map( A1 => n238, A2 => n5014, B1 => n9788, B2 => 
                           n5015, ZN => n9841);
   U10983 : NAND3_X1 port map( A1 => n9845, A2 => n9846, A3 => n9847, ZN => 
                           n12145);
   U10984 : AOI221_X1 port map( B1 => n9783, B2 => n5019, C1 => n174, C2 => 
                           MEM_IN(15), A => n9848, ZN => n9847);
   U10985 : OAI22_X1 port map( A1 => n10782, A2 => n257, B1 => n5021, B2 => 
                           n129, ZN => n9848);
   U10986 : AOI22_X1 port map( A1 => n9786, A2 => n5022, B1 => n9787, B2 => 
                           n5023, ZN => n9846);
   U10987 : AOI22_X1 port map( A1 => n238, A2 => n5024, B1 => n9788, B2 => 
                           n5025, ZN => n9845);
   U10988 : NAND3_X1 port map( A1 => n9849, A2 => n9850, A3 => n9851, ZN => 
                           n12144);
   U10989 : AOI221_X1 port map( B1 => n9783, B2 => n5029, C1 => n174, C2 => 
                           MEM_IN(16), A => n9852, ZN => n9851);
   U10990 : OAI22_X1 port map( A1 => n10781, A2 => n257, B1 => n5031, B2 => 
                           n129, ZN => n9852);
   U10991 : AOI22_X1 port map( A1 => n9786, A2 => n5032, B1 => n9787, B2 => 
                           n5033, ZN => n9850);
   U10992 : AOI22_X1 port map( A1 => n238, A2 => n5034, B1 => n9788, B2 => 
                           n5035, ZN => n9849);
   U10993 : NAND3_X1 port map( A1 => n9853, A2 => n9854, A3 => n9855, ZN => 
                           n12143);
   U10994 : AOI221_X1 port map( B1 => n9783, B2 => n5039, C1 => n174, C2 => 
                           MEM_IN(17), A => n9856, ZN => n9855);
   U10995 : OAI22_X1 port map( A1 => n10780, A2 => n257, B1 => n5041, B2 => 
                           n129, ZN => n9856);
   U10996 : AOI22_X1 port map( A1 => n9786, A2 => n5042, B1 => n9787, B2 => 
                           n5043, ZN => n9854);
   U10997 : AOI22_X1 port map( A1 => n238, A2 => n5044, B1 => n9788, B2 => 
                           n5045, ZN => n9853);
   U10998 : NAND3_X1 port map( A1 => n9857, A2 => n9858, A3 => n9859, ZN => 
                           n12142);
   U10999 : AOI221_X1 port map( B1 => n9783, B2 => n5049, C1 => n174, C2 => 
                           MEM_IN(18), A => n9860, ZN => n9859);
   U11000 : OAI22_X1 port map( A1 => n10779, A2 => n257, B1 => n5051, B2 => 
                           n129, ZN => n9860);
   U11001 : AOI22_X1 port map( A1 => n9786, A2 => n5052, B1 => n9787, B2 => 
                           n5053, ZN => n9858);
   U11002 : AOI22_X1 port map( A1 => n238, A2 => n5054, B1 => n9788, B2 => 
                           n5055, ZN => n9857);
   U11003 : NAND3_X1 port map( A1 => n9861, A2 => n9862, A3 => n9863, ZN => 
                           n12141);
   U11004 : AOI221_X1 port map( B1 => n9783, B2 => n5059, C1 => n174, C2 => 
                           MEM_IN(19), A => n9864, ZN => n9863);
   U11005 : OAI22_X1 port map( A1 => n10778, A2 => n257, B1 => n5061, B2 => 
                           n129, ZN => n9864);
   U11006 : AOI22_X1 port map( A1 => n9786, A2 => n5062, B1 => n9787, B2 => 
                           n5063, ZN => n9862);
   U11007 : AOI22_X1 port map( A1 => n238, A2 => n5064, B1 => n9788, B2 => 
                           n5065, ZN => n9861);
   U11008 : NAND3_X1 port map( A1 => n9865, A2 => n9866, A3 => n9867, ZN => 
                           n12140);
   U11009 : AOI221_X1 port map( B1 => n9783, B2 => n5069, C1 => n174, C2 => 
                           MEM_IN(20), A => n9868, ZN => n9867);
   U11010 : OAI22_X1 port map( A1 => n10777, A2 => n257, B1 => n5071, B2 => 
                           n129, ZN => n9868);
   U11011 : AOI22_X1 port map( A1 => n9786, A2 => n5072, B1 => n9787, B2 => 
                           n5073, ZN => n9866);
   U11012 : AOI22_X1 port map( A1 => n238, A2 => n5074, B1 => n9788, B2 => 
                           n5075, ZN => n9865);
   U11013 : NAND3_X1 port map( A1 => n9869, A2 => n9870, A3 => n9871, ZN => 
                           n12139);
   U11014 : AOI221_X1 port map( B1 => n9783, B2 => n5079, C1 => n174, C2 => 
                           MEM_IN(21), A => n9872, ZN => n9871);
   U11015 : OAI22_X1 port map( A1 => n10776, A2 => n257, B1 => n5081, B2 => 
                           n129, ZN => n9872);
   U11016 : AOI22_X1 port map( A1 => n9786, A2 => n5082, B1 => n9787, B2 => 
                           n5083, ZN => n9870);
   U11017 : AOI22_X1 port map( A1 => n238, A2 => n5084, B1 => n9788, B2 => 
                           n5085, ZN => n9869);
   U11018 : NAND3_X1 port map( A1 => n9873, A2 => n9874, A3 => n9875, ZN => 
                           n12138);
   U11019 : AOI221_X1 port map( B1 => n9783, B2 => n5089, C1 => n174, C2 => 
                           MEM_IN(22), A => n9876, ZN => n9875);
   U11020 : OAI22_X1 port map( A1 => n10775, A2 => n257, B1 => n5091, B2 => 
                           n129, ZN => n9876);
   U11021 : AOI22_X1 port map( A1 => n9786, A2 => n5092, B1 => n9787, B2 => 
                           n5093, ZN => n9874);
   U11022 : AOI22_X1 port map( A1 => n238, A2 => n5094, B1 => n9788, B2 => 
                           n5095, ZN => n9873);
   U11023 : NAND3_X1 port map( A1 => n9877, A2 => n9878, A3 => n9879, ZN => 
                           n12137);
   U11024 : AOI221_X1 port map( B1 => n9783, B2 => n5099, C1 => n174, C2 => 
                           MEM_IN(23), A => n9880, ZN => n9879);
   U11025 : OAI22_X1 port map( A1 => n10774, A2 => n257, B1 => n5101, B2 => 
                           n129, ZN => n9880);
   U11026 : AOI22_X1 port map( A1 => n9786, A2 => n5102, B1 => n9787, B2 => 
                           n5103, ZN => n9878);
   U11027 : AOI22_X1 port map( A1 => n238, A2 => n5104, B1 => n9788, B2 => 
                           n5105, ZN => n9877);
   U11028 : NAND3_X1 port map( A1 => n9881, A2 => n9882, A3 => n9883, ZN => 
                           n12136);
   U11029 : AOI221_X1 port map( B1 => n9783, B2 => n5109, C1 => n174, C2 => 
                           MEM_IN(24), A => n9884, ZN => n9883);
   U11030 : OAI22_X1 port map( A1 => n10773, A2 => n257, B1 => n5111, B2 => 
                           n129, ZN => n9884);
   U11031 : AOI22_X1 port map( A1 => n9786, A2 => n5112, B1 => n9787, B2 => 
                           n5113, ZN => n9882);
   U11032 : AOI22_X1 port map( A1 => n238, A2 => n5114, B1 => n9788, B2 => 
                           n5115, ZN => n9881);
   U11033 : NAND3_X1 port map( A1 => n9885, A2 => n9886, A3 => n9887, ZN => 
                           n12135);
   U11034 : AOI221_X1 port map( B1 => n9783, B2 => n5119, C1 => n174, C2 => 
                           MEM_IN(25), A => n9888, ZN => n9887);
   U11035 : OAI22_X1 port map( A1 => n10772, A2 => n257, B1 => n5121, B2 => 
                           n129, ZN => n9888);
   U11036 : AOI22_X1 port map( A1 => n9786, A2 => n5122, B1 => n9787, B2 => 
                           n5123, ZN => n9886);
   U11037 : AOI22_X1 port map( A1 => n238, A2 => n5124, B1 => n9788, B2 => 
                           n5125, ZN => n9885);
   U11038 : NAND3_X1 port map( A1 => n9889, A2 => n9890, A3 => n9891, ZN => 
                           n12134);
   U11039 : AOI221_X1 port map( B1 => n9783, B2 => n5129, C1 => n174, C2 => 
                           MEM_IN(26), A => n9892, ZN => n9891);
   U11040 : OAI22_X1 port map( A1 => n10771, A2 => n257, B1 => n5131, B2 => 
                           n129, ZN => n9892);
   U11041 : AOI22_X1 port map( A1 => n9786, A2 => n5132, B1 => n9787, B2 => 
                           n5133, ZN => n9890);
   U11042 : AOI22_X1 port map( A1 => n238, A2 => n5134, B1 => n9788, B2 => 
                           n5135, ZN => n9889);
   U11043 : NAND3_X1 port map( A1 => n9893, A2 => n9894, A3 => n9895, ZN => 
                           n12133);
   U11044 : AOI221_X1 port map( B1 => n9783, B2 => n5139, C1 => n174, C2 => 
                           MEM_IN(27), A => n9896, ZN => n9895);
   U11045 : OAI22_X1 port map( A1 => n10770, A2 => n257, B1 => n5141, B2 => 
                           n129, ZN => n9896);
   U11046 : AOI22_X1 port map( A1 => n9786, A2 => n5142, B1 => n9787, B2 => 
                           n5143, ZN => n9894);
   U11047 : AOI22_X1 port map( A1 => n238, A2 => n5144, B1 => n9788, B2 => 
                           n5145, ZN => n9893);
   U11048 : NAND3_X1 port map( A1 => n9897, A2 => n9898, A3 => n9899, ZN => 
                           n12132);
   U11049 : AOI221_X1 port map( B1 => n9783, B2 => n5149, C1 => n174, C2 => 
                           MEM_IN(28), A => n9900, ZN => n9899);
   U11050 : OAI22_X1 port map( A1 => n10769, A2 => n257, B1 => n5151, B2 => 
                           n129, ZN => n9900);
   U11051 : AOI22_X1 port map( A1 => n9786, A2 => n5152, B1 => n9787, B2 => 
                           n5153, ZN => n9898);
   U11052 : AOI22_X1 port map( A1 => n238, A2 => n5154, B1 => n9788, B2 => 
                           n5155, ZN => n9897);
   U11053 : NAND3_X1 port map( A1 => n9901, A2 => n9902, A3 => n9903, ZN => 
                           n12131);
   U11054 : AOI221_X1 port map( B1 => n9783, B2 => n5159, C1 => n174, C2 => 
                           MEM_IN(29), A => n9904, ZN => n9903);
   U11055 : OAI22_X1 port map( A1 => n10768, A2 => n257, B1 => n5161, B2 => 
                           n129, ZN => n9904);
   U11056 : AOI22_X1 port map( A1 => n9786, A2 => n5162, B1 => n9787, B2 => 
                           n5163, ZN => n9902);
   U11057 : AOI22_X1 port map( A1 => n238, A2 => n5164, B1 => n9788, B2 => 
                           n5165, ZN => n9901);
   U11058 : NAND3_X1 port map( A1 => n9905, A2 => n9906, A3 => n9907, ZN => 
                           n12130);
   U11059 : AOI221_X1 port map( B1 => n9783, B2 => n5169, C1 => n174, C2 => 
                           MEM_IN(30), A => n9908, ZN => n9907);
   U11060 : OAI22_X1 port map( A1 => n10767, A2 => n257, B1 => n5171, B2 => 
                           n129, ZN => n9908);
   U11061 : AOI22_X1 port map( A1 => n9786, A2 => n5172, B1 => n9787, B2 => 
                           n5173, ZN => n9906);
   U11062 : AOI22_X1 port map( A1 => n238, A2 => n5174, B1 => n9788, B2 => 
                           n5175, ZN => n9905);
   U11063 : NAND3_X1 port map( A1 => n9909, A2 => n9910, A3 => n9911, ZN => 
                           n12129);
   U11064 : AOI221_X1 port map( B1 => n9783, B2 => n5179, C1 => n174, C2 => 
                           MEM_IN(31), A => n9912, ZN => n9911);
   U11065 : OAI22_X1 port map( A1 => n10766, A2 => n257, B1 => n5181, B2 => 
                           n129, ZN => n9912);
   U11066 : AOI22_X1 port map( A1 => n9786, A2 => n5191, B1 => n9787, B2 => 
                           n5192, ZN => n9910);
   U11067 : AOI22_X1 port map( A1 => n238, A2 => n5195, B1 => n9788, B2 => 
                           n5196, ZN => n9909);
   U11068 : INV_X1 port map( A => n9920, ZN => n9917);
   U11069 : AOI22_X1 port map( A1 => n9915, A2 => n9922, B1 => n4841, B2 => 
                           n257, ZN => n9920);
   U11070 : INV_X1 port map( A => n9914, ZN => n9922);
   U11071 : NAND3_X1 port map( A1 => n208, A2 => n257, A3 => n8893, ZN => n9914
                           );
   U11072 : INV_X1 port map( A => n9913, ZN => n8893);
   U11073 : OAI22_X1 port map( A1 => n9923, A2 => n4786, B1 => n9924, B2 => 
                           n5204, ZN => n9785);
   U11074 : NOR2_X1 port map( A1 => n9913, A2 => n9925, ZN => n9924);
   U11075 : INV_X1 port map( A => n9915, ZN => n9925);
   U11076 : NAND4_X1 port map( A1 => n9775, A2 => n9779, A3 => n9192, A4 => 
                           n9045, ZN => n9913);
   U11077 : NOR4_X1 port map( A1 => n9926, A2 => n9772, A3 => RESET, A4 => 
                           n9918, ZN => n9923);
   U11078 : OAI211_X1 port map( C1 => n6374, C2 => n9043, A => n9475, B => 
                           n9623, ZN => n9926);
   U11079 : INV_X1 port map( A => n9482, ZN => n9475);
   U11080 : NOR2_X1 port map( A1 => n9045, A2 => n4787, ZN => n9482);
   U11081 : NAND3_X1 port map( A1 => n6377, A2 => n8743, A3 => n7560, ZN => 
                           n9043);
   U11082 : INV_X1 port map( A => n8742, ZN => n6377);
   U11083 : NOR2_X1 port map( A1 => n9927, A2 => n9928, ZN => n9915);
   U11084 : NAND2_X1 port map( A1 => n8895, A2 => n6381, ZN => n9045);
   U11085 : NAND3_X1 port map( A1 => n9929, A2 => n9930, A3 => n9931, ZN => 
                           n12128);
   U11086 : AOI221_X1 port map( B1 => n9932, B2 => n4863, C1 => n175, C2 => 
                           MEM_IN(0), A => n9933, ZN => n9931);
   U11087 : OAI22_X1 port map( A1 => n10765, A2 => n271, B1 => n4867, B2 => 
                           n126, ZN => n9933);
   U11088 : AOI22_X1 port map( A1 => n9935, A2 => n4869, B1 => n9936, B2 => 
                           n4871, ZN => n9930);
   U11089 : AOI22_X1 port map( A1 => n9937, A2 => n4873, B1 => n9938, B2 => 
                           n4875, ZN => n9929);
   U11090 : NAND3_X1 port map( A1 => n9939, A2 => n9940, A3 => n9941, ZN => 
                           n12127);
   U11091 : AOI221_X1 port map( B1 => n9932, B2 => n4879, C1 => n175, C2 => 
                           MEM_IN(1), A => n9942, ZN => n9941);
   U11092 : OAI22_X1 port map( A1 => n10764, A2 => n271, B1 => n4881, B2 => 
                           n126, ZN => n9942);
   U11093 : AOI22_X1 port map( A1 => n9935, A2 => n4882, B1 => n9936, B2 => 
                           n4883, ZN => n9940);
   U11094 : AOI22_X1 port map( A1 => n9937, A2 => n4884, B1 => n9938, B2 => 
                           n4885, ZN => n9939);
   U11095 : NAND3_X1 port map( A1 => n9943, A2 => n9944, A3 => n9945, ZN => 
                           n12126);
   U11096 : AOI221_X1 port map( B1 => n9932, B2 => n4889, C1 => n175, C2 => 
                           MEM_IN(2), A => n9946, ZN => n9945);
   U11097 : OAI22_X1 port map( A1 => n10763, A2 => n271, B1 => n4891, B2 => 
                           n126, ZN => n9946);
   U11098 : AOI22_X1 port map( A1 => n9935, A2 => n4892, B1 => n9936, B2 => 
                           n4893, ZN => n9944);
   U11099 : AOI22_X1 port map( A1 => n9937, A2 => n4894, B1 => n9938, B2 => 
                           n4895, ZN => n9943);
   U11100 : NAND3_X1 port map( A1 => n9947, A2 => n9948, A3 => n9949, ZN => 
                           n12125);
   U11101 : AOI221_X1 port map( B1 => n9932, B2 => n4899, C1 => n175, C2 => 
                           MEM_IN(3), A => n9950, ZN => n9949);
   U11102 : OAI22_X1 port map( A1 => n10762, A2 => n271, B1 => n4901, B2 => 
                           n126, ZN => n9950);
   U11103 : AOI22_X1 port map( A1 => n9935, A2 => n4902, B1 => n9936, B2 => 
                           n4903, ZN => n9948);
   U11104 : AOI22_X1 port map( A1 => n9937, A2 => n4904, B1 => n9938, B2 => 
                           n4905, ZN => n9947);
   U11105 : NAND3_X1 port map( A1 => n9951, A2 => n9952, A3 => n9953, ZN => 
                           n12124);
   U11106 : AOI221_X1 port map( B1 => n9932, B2 => n4909, C1 => n175, C2 => 
                           MEM_IN(4), A => n9954, ZN => n9953);
   U11107 : OAI22_X1 port map( A1 => n10761, A2 => n271, B1 => n4911, B2 => 
                           n126, ZN => n9954);
   U11108 : AOI22_X1 port map( A1 => n9935, A2 => n4912, B1 => n9936, B2 => 
                           n4913, ZN => n9952);
   U11109 : AOI22_X1 port map( A1 => n9937, A2 => n4914, B1 => n9938, B2 => 
                           n4915, ZN => n9951);
   U11110 : NAND3_X1 port map( A1 => n9955, A2 => n9956, A3 => n9957, ZN => 
                           n12123);
   U11111 : AOI221_X1 port map( B1 => n9932, B2 => n4919, C1 => n175, C2 => 
                           MEM_IN(5), A => n9958, ZN => n9957);
   U11112 : OAI22_X1 port map( A1 => n10760, A2 => n271, B1 => n4921, B2 => 
                           n126, ZN => n9958);
   U11113 : AOI22_X1 port map( A1 => n9935, A2 => n4922, B1 => n9936, B2 => 
                           n4923, ZN => n9956);
   U11114 : AOI22_X1 port map( A1 => n9937, A2 => n4924, B1 => n9938, B2 => 
                           n4925, ZN => n9955);
   U11115 : NAND3_X1 port map( A1 => n9959, A2 => n9960, A3 => n9961, ZN => 
                           n12122);
   U11116 : AOI221_X1 port map( B1 => n9932, B2 => n4929, C1 => n175, C2 => 
                           MEM_IN(6), A => n9962, ZN => n9961);
   U11117 : OAI22_X1 port map( A1 => n10759, A2 => n271, B1 => n4931, B2 => 
                           n126, ZN => n9962);
   U11118 : AOI22_X1 port map( A1 => n9935, A2 => n4932, B1 => n9936, B2 => 
                           n4933, ZN => n9960);
   U11119 : AOI22_X1 port map( A1 => n9937, A2 => n4934, B1 => n9938, B2 => 
                           n4935, ZN => n9959);
   U11120 : NAND3_X1 port map( A1 => n9963, A2 => n9964, A3 => n9965, ZN => 
                           n12121);
   U11121 : AOI221_X1 port map( B1 => n9932, B2 => n4939, C1 => n175, C2 => 
                           MEM_IN(7), A => n9966, ZN => n9965);
   U11122 : OAI22_X1 port map( A1 => n10758, A2 => n271, B1 => n4941, B2 => 
                           n126, ZN => n9966);
   U11123 : AOI22_X1 port map( A1 => n9935, A2 => n4942, B1 => n9936, B2 => 
                           n4943, ZN => n9964);
   U11124 : AOI22_X1 port map( A1 => n9937, A2 => n4944, B1 => n9938, B2 => 
                           n4945, ZN => n9963);
   U11125 : NAND3_X1 port map( A1 => n9967, A2 => n9968, A3 => n9969, ZN => 
                           n12120);
   U11126 : AOI221_X1 port map( B1 => n9932, B2 => n4949, C1 => n175, C2 => 
                           MEM_IN(8), A => n9970, ZN => n9969);
   U11127 : OAI22_X1 port map( A1 => n10757, A2 => n271, B1 => n4951, B2 => 
                           n126, ZN => n9970);
   U11128 : AOI22_X1 port map( A1 => n9935, A2 => n4952, B1 => n9936, B2 => 
                           n4953, ZN => n9968);
   U11129 : AOI22_X1 port map( A1 => n9937, A2 => n4954, B1 => n9938, B2 => 
                           n4955, ZN => n9967);
   U11130 : NAND3_X1 port map( A1 => n9971, A2 => n9972, A3 => n9973, ZN => 
                           n12119);
   U11131 : AOI221_X1 port map( B1 => n9932, B2 => n4959, C1 => n175, C2 => 
                           MEM_IN(9), A => n9974, ZN => n9973);
   U11132 : OAI22_X1 port map( A1 => n10756, A2 => n271, B1 => n4961, B2 => 
                           n126, ZN => n9974);
   U11133 : AOI22_X1 port map( A1 => n9935, A2 => n4962, B1 => n9936, B2 => 
                           n4963, ZN => n9972);
   U11134 : AOI22_X1 port map( A1 => n9937, A2 => n4964, B1 => n9938, B2 => 
                           n4965, ZN => n9971);
   U11135 : NAND3_X1 port map( A1 => n9975, A2 => n9976, A3 => n9977, ZN => 
                           n12118);
   U11136 : AOI221_X1 port map( B1 => n9932, B2 => n4969, C1 => n175, C2 => 
                           MEM_IN(10), A => n9978, ZN => n9977);
   U11137 : OAI22_X1 port map( A1 => n10755, A2 => n271, B1 => n4971, B2 => 
                           n126, ZN => n9978);
   U11138 : AOI22_X1 port map( A1 => n9935, A2 => n4972, B1 => n9936, B2 => 
                           n4973, ZN => n9976);
   U11139 : AOI22_X1 port map( A1 => n9937, A2 => n4974, B1 => n9938, B2 => 
                           n4975, ZN => n9975);
   U11140 : NAND3_X1 port map( A1 => n9979, A2 => n9980, A3 => n9981, ZN => 
                           n12117);
   U11141 : AOI221_X1 port map( B1 => n9932, B2 => n4979, C1 => n175, C2 => 
                           MEM_IN(11), A => n9982, ZN => n9981);
   U11142 : OAI22_X1 port map( A1 => n10754, A2 => n271, B1 => n4981, B2 => 
                           n126, ZN => n9982);
   U11143 : AOI22_X1 port map( A1 => n9935, A2 => n4982, B1 => n9936, B2 => 
                           n4983, ZN => n9980);
   U11144 : AOI22_X1 port map( A1 => n9937, A2 => n4984, B1 => n9938, B2 => 
                           n4985, ZN => n9979);
   U11145 : NAND3_X1 port map( A1 => n9983, A2 => n9984, A3 => n9985, ZN => 
                           n12116);
   U11146 : AOI221_X1 port map( B1 => n9932, B2 => n4989, C1 => n175, C2 => 
                           MEM_IN(12), A => n9986, ZN => n9985);
   U11147 : OAI22_X1 port map( A1 => n10753, A2 => n271, B1 => n4991, B2 => 
                           n126, ZN => n9986);
   U11148 : AOI22_X1 port map( A1 => n9935, A2 => n4992, B1 => n9936, B2 => 
                           n4993, ZN => n9984);
   U11149 : AOI22_X1 port map( A1 => n9937, A2 => n4994, B1 => n9938, B2 => 
                           n4995, ZN => n9983);
   U11150 : NAND3_X1 port map( A1 => n9987, A2 => n9988, A3 => n9989, ZN => 
                           n12115);
   U11151 : AOI221_X1 port map( B1 => n9932, B2 => n4999, C1 => n175, C2 => 
                           MEM_IN(13), A => n9990, ZN => n9989);
   U11152 : OAI22_X1 port map( A1 => n10752, A2 => n271, B1 => n5001, B2 => 
                           n126, ZN => n9990);
   U11153 : AOI22_X1 port map( A1 => n9935, A2 => n5002, B1 => n9936, B2 => 
                           n5003, ZN => n9988);
   U11154 : AOI22_X1 port map( A1 => n9937, A2 => n5004, B1 => n9938, B2 => 
                           n5005, ZN => n9987);
   U11155 : NAND3_X1 port map( A1 => n9991, A2 => n9992, A3 => n9993, ZN => 
                           n12114);
   U11156 : AOI221_X1 port map( B1 => n9932, B2 => n5009, C1 => n175, C2 => 
                           MEM_IN(14), A => n9994, ZN => n9993);
   U11157 : OAI22_X1 port map( A1 => n10751, A2 => n271, B1 => n5011, B2 => 
                           n126, ZN => n9994);
   U11158 : AOI22_X1 port map( A1 => n9935, A2 => n5012, B1 => n9936, B2 => 
                           n5013, ZN => n9992);
   U11159 : AOI22_X1 port map( A1 => n9937, A2 => n5014, B1 => n9938, B2 => 
                           n5015, ZN => n9991);
   U11160 : NAND3_X1 port map( A1 => n9995, A2 => n9996, A3 => n9997, ZN => 
                           n12113);
   U11161 : AOI221_X1 port map( B1 => n9932, B2 => n5019, C1 => n175, C2 => 
                           MEM_IN(15), A => n9998, ZN => n9997);
   U11162 : OAI22_X1 port map( A1 => n10750, A2 => n271, B1 => n5021, B2 => 
                           n126, ZN => n9998);
   U11163 : AOI22_X1 port map( A1 => n9935, A2 => n5022, B1 => n9936, B2 => 
                           n5023, ZN => n9996);
   U11164 : AOI22_X1 port map( A1 => n9937, A2 => n5024, B1 => n9938, B2 => 
                           n5025, ZN => n9995);
   U11165 : NAND3_X1 port map( A1 => n9999, A2 => n10000, A3 => n10001, ZN => 
                           n12112);
   U11166 : AOI221_X1 port map( B1 => n9932, B2 => n5029, C1 => n175, C2 => 
                           MEM_IN(16), A => n10002, ZN => n10001);
   U11167 : OAI22_X1 port map( A1 => n10749, A2 => n271, B1 => n5031, B2 => 
                           n126, ZN => n10002);
   U11168 : AOI22_X1 port map( A1 => n9935, A2 => n5032, B1 => n9936, B2 => 
                           n5033, ZN => n10000);
   U11169 : AOI22_X1 port map( A1 => n9937, A2 => n5034, B1 => n9938, B2 => 
                           n5035, ZN => n9999);
   U11170 : NAND3_X1 port map( A1 => n10003, A2 => n10004, A3 => n10005, ZN => 
                           n12111);
   U11171 : AOI221_X1 port map( B1 => n9932, B2 => n5039, C1 => n175, C2 => 
                           MEM_IN(17), A => n10006, ZN => n10005);
   U11172 : OAI22_X1 port map( A1 => n10748, A2 => n271, B1 => n5041, B2 => 
                           n126, ZN => n10006);
   U11173 : AOI22_X1 port map( A1 => n9935, A2 => n5042, B1 => n9936, B2 => 
                           n5043, ZN => n10004);
   U11174 : AOI22_X1 port map( A1 => n9937, A2 => n5044, B1 => n9938, B2 => 
                           n5045, ZN => n10003);
   U11175 : NAND3_X1 port map( A1 => n10007, A2 => n10008, A3 => n10009, ZN => 
                           n12110);
   U11176 : AOI221_X1 port map( B1 => n9932, B2 => n5049, C1 => n175, C2 => 
                           MEM_IN(18), A => n10010, ZN => n10009);
   U11177 : OAI22_X1 port map( A1 => n10747, A2 => n271, B1 => n5051, B2 => 
                           n126, ZN => n10010);
   U11178 : AOI22_X1 port map( A1 => n9935, A2 => n5052, B1 => n9936, B2 => 
                           n5053, ZN => n10008);
   U11179 : AOI22_X1 port map( A1 => n9937, A2 => n5054, B1 => n9938, B2 => 
                           n5055, ZN => n10007);
   U11180 : NAND3_X1 port map( A1 => n10011, A2 => n10012, A3 => n10013, ZN => 
                           n12109);
   U11181 : AOI221_X1 port map( B1 => n9932, B2 => n5059, C1 => n175, C2 => 
                           MEM_IN(19), A => n10014, ZN => n10013);
   U11182 : OAI22_X1 port map( A1 => n10746, A2 => n271, B1 => n5061, B2 => 
                           n126, ZN => n10014);
   U11183 : AOI22_X1 port map( A1 => n9935, A2 => n5062, B1 => n9936, B2 => 
                           n5063, ZN => n10012);
   U11184 : AOI22_X1 port map( A1 => n9937, A2 => n5064, B1 => n9938, B2 => 
                           n5065, ZN => n10011);
   U11185 : NAND3_X1 port map( A1 => n10015, A2 => n10016, A3 => n10017, ZN => 
                           n12108);
   U11186 : AOI221_X1 port map( B1 => n9932, B2 => n5069, C1 => n175, C2 => 
                           MEM_IN(20), A => n10018, ZN => n10017);
   U11187 : OAI22_X1 port map( A1 => n10745, A2 => n271, B1 => n5071, B2 => 
                           n126, ZN => n10018);
   U11188 : AOI22_X1 port map( A1 => n9935, A2 => n5072, B1 => n9936, B2 => 
                           n5073, ZN => n10016);
   U11189 : AOI22_X1 port map( A1 => n9937, A2 => n5074, B1 => n9938, B2 => 
                           n5075, ZN => n10015);
   U11190 : NAND3_X1 port map( A1 => n10019, A2 => n10020, A3 => n10021, ZN => 
                           n12107);
   U11191 : AOI221_X1 port map( B1 => n9932, B2 => n5079, C1 => n175, C2 => 
                           MEM_IN(21), A => n10022, ZN => n10021);
   U11192 : OAI22_X1 port map( A1 => n10744, A2 => n271, B1 => n5081, B2 => 
                           n126, ZN => n10022);
   U11193 : AOI22_X1 port map( A1 => n9935, A2 => n5082, B1 => n9936, B2 => 
                           n5083, ZN => n10020);
   U11194 : AOI22_X1 port map( A1 => n9937, A2 => n5084, B1 => n9938, B2 => 
                           n5085, ZN => n10019);
   U11195 : NAND3_X1 port map( A1 => n10023, A2 => n10024, A3 => n10025, ZN => 
                           n12106);
   U11196 : AOI221_X1 port map( B1 => n9932, B2 => n5089, C1 => n175, C2 => 
                           MEM_IN(22), A => n10026, ZN => n10025);
   U11197 : OAI22_X1 port map( A1 => n10743, A2 => n271, B1 => n5091, B2 => 
                           n126, ZN => n10026);
   U11198 : AOI22_X1 port map( A1 => n9935, A2 => n5092, B1 => n9936, B2 => 
                           n5093, ZN => n10024);
   U11199 : AOI22_X1 port map( A1 => n9937, A2 => n5094, B1 => n9938, B2 => 
                           n5095, ZN => n10023);
   U11200 : NAND3_X1 port map( A1 => n10027, A2 => n10028, A3 => n10029, ZN => 
                           n12105);
   U11201 : AOI221_X1 port map( B1 => n9932, B2 => n5099, C1 => n175, C2 => 
                           MEM_IN(23), A => n10030, ZN => n10029);
   U11202 : OAI22_X1 port map( A1 => n10742, A2 => n271, B1 => n5101, B2 => 
                           n126, ZN => n10030);
   U11203 : AOI22_X1 port map( A1 => n9935, A2 => n5102, B1 => n9936, B2 => 
                           n5103, ZN => n10028);
   U11204 : AOI22_X1 port map( A1 => n9937, A2 => n5104, B1 => n9938, B2 => 
                           n5105, ZN => n10027);
   U11205 : NAND3_X1 port map( A1 => n10031, A2 => n10032, A3 => n10033, ZN => 
                           n12104);
   U11206 : AOI221_X1 port map( B1 => n9932, B2 => n5109, C1 => n175, C2 => 
                           MEM_IN(24), A => n10034, ZN => n10033);
   U11207 : OAI22_X1 port map( A1 => n10741, A2 => n271, B1 => n5111, B2 => 
                           n126, ZN => n10034);
   U11208 : AOI22_X1 port map( A1 => n9935, A2 => n5112, B1 => n9936, B2 => 
                           n5113, ZN => n10032);
   U11209 : AOI22_X1 port map( A1 => n9937, A2 => n5114, B1 => n9938, B2 => 
                           n5115, ZN => n10031);
   U11210 : NAND3_X1 port map( A1 => n10035, A2 => n10036, A3 => n10037, ZN => 
                           n12103);
   U11211 : AOI221_X1 port map( B1 => n9932, B2 => n5119, C1 => n175, C2 => 
                           MEM_IN(25), A => n10038, ZN => n10037);
   U11212 : OAI22_X1 port map( A1 => n10740, A2 => n271, B1 => n5121, B2 => 
                           n126, ZN => n10038);
   U11213 : AOI22_X1 port map( A1 => n9935, A2 => n5122, B1 => n9936, B2 => 
                           n5123, ZN => n10036);
   U11214 : AOI22_X1 port map( A1 => n9937, A2 => n5124, B1 => n9938, B2 => 
                           n5125, ZN => n10035);
   U11215 : NAND3_X1 port map( A1 => n10039, A2 => n10040, A3 => n10041, ZN => 
                           n12102);
   U11216 : AOI221_X1 port map( B1 => n9932, B2 => n5129, C1 => n175, C2 => 
                           MEM_IN(26), A => n10042, ZN => n10041);
   U11217 : OAI22_X1 port map( A1 => n10739, A2 => n271, B1 => n5131, B2 => 
                           n126, ZN => n10042);
   U11218 : AOI22_X1 port map( A1 => n9935, A2 => n5132, B1 => n9936, B2 => 
                           n5133, ZN => n10040);
   U11219 : AOI22_X1 port map( A1 => n9937, A2 => n5134, B1 => n9938, B2 => 
                           n5135, ZN => n10039);
   U11220 : NAND3_X1 port map( A1 => n10043, A2 => n10044, A3 => n10045, ZN => 
                           n12101);
   U11221 : AOI221_X1 port map( B1 => n9932, B2 => n5139, C1 => n175, C2 => 
                           MEM_IN(27), A => n10046, ZN => n10045);
   U11222 : OAI22_X1 port map( A1 => n10738, A2 => n271, B1 => n5141, B2 => 
                           n126, ZN => n10046);
   U11223 : AOI22_X1 port map( A1 => n9935, A2 => n5142, B1 => n9936, B2 => 
                           n5143, ZN => n10044);
   U11224 : AOI22_X1 port map( A1 => n9937, A2 => n5144, B1 => n9938, B2 => 
                           n5145, ZN => n10043);
   U11225 : NAND3_X1 port map( A1 => n10047, A2 => n10048, A3 => n10049, ZN => 
                           n12100);
   U11226 : AOI221_X1 port map( B1 => n9932, B2 => n5149, C1 => n175, C2 => 
                           MEM_IN(28), A => n10050, ZN => n10049);
   U11227 : OAI22_X1 port map( A1 => n10737, A2 => n271, B1 => n5151, B2 => 
                           n126, ZN => n10050);
   U11228 : AOI22_X1 port map( A1 => n9935, A2 => n5152, B1 => n9936, B2 => 
                           n5153, ZN => n10048);
   U11229 : AOI22_X1 port map( A1 => n9937, A2 => n5154, B1 => n9938, B2 => 
                           n5155, ZN => n10047);
   U11230 : NAND3_X1 port map( A1 => n10051, A2 => n10052, A3 => n10053, ZN => 
                           n12099);
   U11231 : AOI221_X1 port map( B1 => n9932, B2 => n5159, C1 => n175, C2 => 
                           MEM_IN(29), A => n10054, ZN => n10053);
   U11232 : OAI22_X1 port map( A1 => n10736, A2 => n271, B1 => n5161, B2 => 
                           n126, ZN => n10054);
   U11233 : AOI22_X1 port map( A1 => n9935, A2 => n5162, B1 => n9936, B2 => 
                           n5163, ZN => n10052);
   U11234 : AOI22_X1 port map( A1 => n9937, A2 => n5164, B1 => n9938, B2 => 
                           n5165, ZN => n10051);
   U11235 : NAND3_X1 port map( A1 => n10055, A2 => n10056, A3 => n10057, ZN => 
                           n12098);
   U11236 : AOI221_X1 port map( B1 => n9932, B2 => n5169, C1 => n175, C2 => 
                           MEM_IN(30), A => n10058, ZN => n10057);
   U11237 : OAI22_X1 port map( A1 => n10735, A2 => n271, B1 => n5171, B2 => 
                           n126, ZN => n10058);
   U11238 : AOI22_X1 port map( A1 => n9935, A2 => n5172, B1 => n9936, B2 => 
                           n5173, ZN => n10056);
   U11239 : AOI22_X1 port map( A1 => n9937, A2 => n5174, B1 => n9938, B2 => 
                           n5175, ZN => n10055);
   U11240 : NAND3_X1 port map( A1 => n10059, A2 => n10060, A3 => n10061, ZN => 
                           n12097);
   U11241 : AOI221_X1 port map( B1 => n9932, B2 => n5179, C1 => n175, C2 => 
                           MEM_IN(31), A => n10062, ZN => n10061);
   U11242 : OAI22_X1 port map( A1 => n10734, A2 => n271, B1 => n5181, B2 => 
                           n126, ZN => n10062);
   U11243 : INV_X1 port map( A => n9625, ZN => n9623);
   U11244 : AOI22_X1 port map( A1 => n9935, A2 => n5191, B1 => n9936, B2 => 
                           n5192, ZN => n10060);
   U11245 : AOI22_X1 port map( A1 => n9937, A2 => n5195, B1 => n9938, B2 => 
                           n5196, ZN => n10059);
   U11246 : OAI22_X1 port map( A1 => n10069, A2 => n10064, B1 => n208, B2 => 
                           n270, ZN => n10066);
   U11247 : NAND3_X1 port map( A1 => n208, A2 => n271, A3 => n9044, ZN => 
                           n10064);
   U11248 : INV_X1 port map( A => n10063, ZN => n9044);
   U11249 : OAI22_X1 port map( A1 => n4786, A2 => n10070, B1 => n10071, B2 => 
                           n5204, ZN => n9934);
   U11250 : NOR2_X1 port map( A1 => n10063, A2 => n10069, ZN => n10071);
   U11251 : NAND3_X1 port map( A1 => n9775, A2 => n9192, A3 => n10072, ZN => 
                           n10063);
   U11252 : AOI211_X1 port map( C1 => n10073, C2 => n5207, A => n10074, B => 
                           n9625, ZN => n10070);
   U11253 : NOR2_X1 port map( A1 => n9192, A2 => n4787, ZN => n9625);
   U11254 : NOR3_X1 port map( A1 => n10075, A2 => n10076, A3 => n10077, ZN => 
                           n5207);
   U11255 : INV_X1 port map( A => n10065, ZN => n10069);
   U11256 : NOR2_X1 port map( A1 => n10078, A2 => n10079, ZN => n10065);
   U11257 : NOR2_X1 port map( A1 => n9921, A2 => n9192, ZN => n9919);
   U11258 : NAND2_X1 port map( A1 => n10080, A2 => n5215, ZN => n9192);
   U11259 : NAND3_X1 port map( A1 => n10081, A2 => n10082, A3 => n10083, ZN => 
                           n12096);
   U11260 : AOI221_X1 port map( B1 => n10084, B2 => n4863, C1 => n172, C2 => 
                           MEM_IN(0), A => n10085, ZN => n10083);
   U11261 : OAI22_X1 port map( A1 => n10733, A2 => n273, B1 => n4867, B2 => 
                           n127, ZN => n10085);
   U11262 : AOI22_X1 port map( A1 => n10087, A2 => n4869, B1 => n10088, B2 => 
                           n4871, ZN => n10082);
   U11263 : AOI22_X1 port map( A1 => n10089, A2 => n4873, B1 => n10090, B2 => 
                           n4875, ZN => n10081);
   U11264 : NAND3_X1 port map( A1 => n10091, A2 => n10092, A3 => n10093, ZN => 
                           n12095);
   U11265 : AOI221_X1 port map( B1 => n10084, B2 => n4879, C1 => n172, C2 => 
                           MEM_IN(1), A => n10094, ZN => n10093);
   U11266 : OAI22_X1 port map( A1 => n10732, A2 => n273, B1 => n4881, B2 => 
                           n127, ZN => n10094);
   U11267 : AOI22_X1 port map( A1 => n10087, A2 => n4882, B1 => n10088, B2 => 
                           n4883, ZN => n10092);
   U11268 : AOI22_X1 port map( A1 => n10089, A2 => n4884, B1 => n10090, B2 => 
                           n4885, ZN => n10091);
   U11269 : NAND3_X1 port map( A1 => n10095, A2 => n10096, A3 => n10097, ZN => 
                           n12094);
   U11270 : AOI221_X1 port map( B1 => n10084, B2 => n4889, C1 => n172, C2 => 
                           MEM_IN(2), A => n10098, ZN => n10097);
   U11271 : OAI22_X1 port map( A1 => n10731, A2 => n273, B1 => n4891, B2 => 
                           n127, ZN => n10098);
   U11272 : AOI22_X1 port map( A1 => n10087, A2 => n4892, B1 => n10088, B2 => 
                           n4893, ZN => n10096);
   U11273 : AOI22_X1 port map( A1 => n10089, A2 => n4894, B1 => n10090, B2 => 
                           n4895, ZN => n10095);
   U11274 : NAND3_X1 port map( A1 => n10099, A2 => n10100, A3 => n10101, ZN => 
                           n12093);
   U11275 : AOI221_X1 port map( B1 => n10084, B2 => n4899, C1 => n172, C2 => 
                           MEM_IN(3), A => n10102, ZN => n10101);
   U11276 : OAI22_X1 port map( A1 => n10730, A2 => n273, B1 => n4901, B2 => 
                           n127, ZN => n10102);
   U11277 : AOI22_X1 port map( A1 => n10087, A2 => n4902, B1 => n10088, B2 => 
                           n4903, ZN => n10100);
   U11278 : AOI22_X1 port map( A1 => n10089, A2 => n4904, B1 => n10090, B2 => 
                           n4905, ZN => n10099);
   U11279 : NAND3_X1 port map( A1 => n10103, A2 => n10104, A3 => n10105, ZN => 
                           n12092);
   U11280 : AOI221_X1 port map( B1 => n10084, B2 => n4909, C1 => n172, C2 => 
                           MEM_IN(4), A => n10106, ZN => n10105);
   U11281 : OAI22_X1 port map( A1 => n10729, A2 => n273, B1 => n4911, B2 => 
                           n127, ZN => n10106);
   U11282 : AOI22_X1 port map( A1 => n10087, A2 => n4912, B1 => n10088, B2 => 
                           n4913, ZN => n10104);
   U11283 : AOI22_X1 port map( A1 => n10089, A2 => n4914, B1 => n10090, B2 => 
                           n4915, ZN => n10103);
   U11284 : NAND3_X1 port map( A1 => n10107, A2 => n10108, A3 => n10109, ZN => 
                           n12091);
   U11285 : AOI221_X1 port map( B1 => n10084, B2 => n4919, C1 => n172, C2 => 
                           MEM_IN(5), A => n10110, ZN => n10109);
   U11286 : OAI22_X1 port map( A1 => n10728, A2 => n273, B1 => n4921, B2 => 
                           n127, ZN => n10110);
   U11287 : AOI22_X1 port map( A1 => n10087, A2 => n4922, B1 => n10088, B2 => 
                           n4923, ZN => n10108);
   U11288 : AOI22_X1 port map( A1 => n10089, A2 => n4924, B1 => n10090, B2 => 
                           n4925, ZN => n10107);
   U11289 : NAND3_X1 port map( A1 => n10111, A2 => n10112, A3 => n10113, ZN => 
                           n12090);
   U11290 : AOI221_X1 port map( B1 => n10084, B2 => n4929, C1 => n172, C2 => 
                           MEM_IN(6), A => n10114, ZN => n10113);
   U11291 : OAI22_X1 port map( A1 => n10727, A2 => n273, B1 => n4931, B2 => 
                           n127, ZN => n10114);
   U11292 : AOI22_X1 port map( A1 => n10087, A2 => n4932, B1 => n10088, B2 => 
                           n4933, ZN => n10112);
   U11293 : AOI22_X1 port map( A1 => n10089, A2 => n4934, B1 => n10090, B2 => 
                           n4935, ZN => n10111);
   U11294 : NAND3_X1 port map( A1 => n10115, A2 => n10116, A3 => n10117, ZN => 
                           n12089);
   U11295 : AOI221_X1 port map( B1 => n10084, B2 => n4939, C1 => n172, C2 => 
                           MEM_IN(7), A => n10118, ZN => n10117);
   U11296 : OAI22_X1 port map( A1 => n10726, A2 => n273, B1 => n4941, B2 => 
                           n127, ZN => n10118);
   U11297 : AOI22_X1 port map( A1 => n10087, A2 => n4942, B1 => n10088, B2 => 
                           n4943, ZN => n10116);
   U11298 : AOI22_X1 port map( A1 => n10089, A2 => n4944, B1 => n10090, B2 => 
                           n4945, ZN => n10115);
   U11299 : NAND3_X1 port map( A1 => n10119, A2 => n10120, A3 => n10121, ZN => 
                           n12088);
   U11300 : AOI221_X1 port map( B1 => n10084, B2 => n4949, C1 => n172, C2 => 
                           MEM_IN(8), A => n10122, ZN => n10121);
   U11301 : OAI22_X1 port map( A1 => n10725, A2 => n273, B1 => n4951, B2 => 
                           n127, ZN => n10122);
   U11302 : AOI22_X1 port map( A1 => n10087, A2 => n4952, B1 => n10088, B2 => 
                           n4953, ZN => n10120);
   U11303 : AOI22_X1 port map( A1 => n10089, A2 => n4954, B1 => n10090, B2 => 
                           n4955, ZN => n10119);
   U11304 : NAND3_X1 port map( A1 => n10123, A2 => n10124, A3 => n10125, ZN => 
                           n12087);
   U11305 : AOI221_X1 port map( B1 => n10084, B2 => n4959, C1 => n172, C2 => 
                           MEM_IN(9), A => n10126, ZN => n10125);
   U11306 : OAI22_X1 port map( A1 => n10724, A2 => n273, B1 => n4961, B2 => 
                           n127, ZN => n10126);
   U11307 : AOI22_X1 port map( A1 => n10087, A2 => n4962, B1 => n10088, B2 => 
                           n4963, ZN => n10124);
   U11308 : AOI22_X1 port map( A1 => n10089, A2 => n4964, B1 => n10090, B2 => 
                           n4965, ZN => n10123);
   U11309 : NAND3_X1 port map( A1 => n10127, A2 => n10128, A3 => n10129, ZN => 
                           n12086);
   U11310 : AOI221_X1 port map( B1 => n10084, B2 => n4969, C1 => n172, C2 => 
                           MEM_IN(10), A => n10130, ZN => n10129);
   U11311 : OAI22_X1 port map( A1 => n10723, A2 => n273, B1 => n4971, B2 => 
                           n127, ZN => n10130);
   U11312 : AOI22_X1 port map( A1 => n10087, A2 => n4972, B1 => n10088, B2 => 
                           n4973, ZN => n10128);
   U11313 : AOI22_X1 port map( A1 => n10089, A2 => n4974, B1 => n10090, B2 => 
                           n4975, ZN => n10127);
   U11314 : NAND3_X1 port map( A1 => n10131, A2 => n10132, A3 => n10133, ZN => 
                           n12085);
   U11315 : AOI221_X1 port map( B1 => n10084, B2 => n4979, C1 => n172, C2 => 
                           MEM_IN(11), A => n10134, ZN => n10133);
   U11316 : OAI22_X1 port map( A1 => n10722, A2 => n273, B1 => n4981, B2 => 
                           n127, ZN => n10134);
   U11317 : AOI22_X1 port map( A1 => n10087, A2 => n4982, B1 => n10088, B2 => 
                           n4983, ZN => n10132);
   U11318 : AOI22_X1 port map( A1 => n10089, A2 => n4984, B1 => n10090, B2 => 
                           n4985, ZN => n10131);
   U11319 : NAND3_X1 port map( A1 => n10135, A2 => n10136, A3 => n10137, ZN => 
                           n12084);
   U11320 : AOI221_X1 port map( B1 => n10084, B2 => n4989, C1 => n172, C2 => 
                           MEM_IN(12), A => n10138, ZN => n10137);
   U11321 : OAI22_X1 port map( A1 => n10721, A2 => n273, B1 => n4991, B2 => 
                           n127, ZN => n10138);
   U11322 : AOI22_X1 port map( A1 => n10087, A2 => n4992, B1 => n10088, B2 => 
                           n4993, ZN => n10136);
   U11323 : AOI22_X1 port map( A1 => n10089, A2 => n4994, B1 => n10090, B2 => 
                           n4995, ZN => n10135);
   U11324 : NAND3_X1 port map( A1 => n10139, A2 => n10140, A3 => n10141, ZN => 
                           n12083);
   U11325 : AOI221_X1 port map( B1 => n10084, B2 => n4999, C1 => n172, C2 => 
                           MEM_IN(13), A => n10142, ZN => n10141);
   U11326 : OAI22_X1 port map( A1 => n10720, A2 => n273, B1 => n5001, B2 => 
                           n127, ZN => n10142);
   U11327 : AOI22_X1 port map( A1 => n10087, A2 => n5002, B1 => n10088, B2 => 
                           n5003, ZN => n10140);
   U11328 : AOI22_X1 port map( A1 => n10089, A2 => n5004, B1 => n10090, B2 => 
                           n5005, ZN => n10139);
   U11329 : NAND3_X1 port map( A1 => n10143, A2 => n10144, A3 => n10145, ZN => 
                           n12082);
   U11330 : AOI221_X1 port map( B1 => n10084, B2 => n5009, C1 => n172, C2 => 
                           MEM_IN(14), A => n10146, ZN => n10145);
   U11331 : OAI22_X1 port map( A1 => n10719, A2 => n273, B1 => n5011, B2 => 
                           n127, ZN => n10146);
   U11332 : AOI22_X1 port map( A1 => n10087, A2 => n5012, B1 => n10088, B2 => 
                           n5013, ZN => n10144);
   U11333 : AOI22_X1 port map( A1 => n10089, A2 => n5014, B1 => n10090, B2 => 
                           n5015, ZN => n10143);
   U11334 : NAND3_X1 port map( A1 => n10147, A2 => n10148, A3 => n10149, ZN => 
                           n12081);
   U11335 : AOI221_X1 port map( B1 => n10084, B2 => n5019, C1 => n172, C2 => 
                           MEM_IN(15), A => n10150, ZN => n10149);
   U11336 : OAI22_X1 port map( A1 => n10718, A2 => n273, B1 => n5021, B2 => 
                           n127, ZN => n10150);
   U11337 : AOI22_X1 port map( A1 => n10087, A2 => n5022, B1 => n10088, B2 => 
                           n5023, ZN => n10148);
   U11338 : AOI22_X1 port map( A1 => n10089, A2 => n5024, B1 => n10090, B2 => 
                           n5025, ZN => n10147);
   U11339 : NAND3_X1 port map( A1 => n10151, A2 => n10152, A3 => n10153, ZN => 
                           n12080);
   U11340 : AOI221_X1 port map( B1 => n10084, B2 => n5029, C1 => n172, C2 => 
                           MEM_IN(16), A => n10154, ZN => n10153);
   U11341 : OAI22_X1 port map( A1 => n10717, A2 => n273, B1 => n5031, B2 => 
                           n127, ZN => n10154);
   U11342 : AOI22_X1 port map( A1 => n10087, A2 => n5032, B1 => n10088, B2 => 
                           n5033, ZN => n10152);
   U11343 : AOI22_X1 port map( A1 => n10089, A2 => n5034, B1 => n10090, B2 => 
                           n5035, ZN => n10151);
   U11344 : NAND3_X1 port map( A1 => n10155, A2 => n10156, A3 => n10157, ZN => 
                           n12079);
   U11345 : AOI221_X1 port map( B1 => n10084, B2 => n5039, C1 => n172, C2 => 
                           MEM_IN(17), A => n10158, ZN => n10157);
   U11346 : OAI22_X1 port map( A1 => n10716, A2 => n273, B1 => n5041, B2 => 
                           n127, ZN => n10158);
   U11347 : AOI22_X1 port map( A1 => n10087, A2 => n5042, B1 => n10088, B2 => 
                           n5043, ZN => n10156);
   U11348 : AOI22_X1 port map( A1 => n10089, A2 => n5044, B1 => n10090, B2 => 
                           n5045, ZN => n10155);
   U11349 : NAND3_X1 port map( A1 => n10159, A2 => n10160, A3 => n10161, ZN => 
                           n12078);
   U11350 : AOI221_X1 port map( B1 => n10084, B2 => n5049, C1 => n172, C2 => 
                           MEM_IN(18), A => n10162, ZN => n10161);
   U11351 : OAI22_X1 port map( A1 => n10715, A2 => n273, B1 => n5051, B2 => 
                           n127, ZN => n10162);
   U11352 : AOI22_X1 port map( A1 => n10087, A2 => n5052, B1 => n10088, B2 => 
                           n5053, ZN => n10160);
   U11353 : AOI22_X1 port map( A1 => n10089, A2 => n5054, B1 => n10090, B2 => 
                           n5055, ZN => n10159);
   U11354 : NAND3_X1 port map( A1 => n10163, A2 => n10164, A3 => n10165, ZN => 
                           n12077);
   U11355 : AOI221_X1 port map( B1 => n10084, B2 => n5059, C1 => n172, C2 => 
                           MEM_IN(19), A => n10166, ZN => n10165);
   U11356 : OAI22_X1 port map( A1 => n10714, A2 => n273, B1 => n5061, B2 => 
                           n127, ZN => n10166);
   U11357 : AOI22_X1 port map( A1 => n10087, A2 => n5062, B1 => n10088, B2 => 
                           n5063, ZN => n10164);
   U11358 : AOI22_X1 port map( A1 => n10089, A2 => n5064, B1 => n10090, B2 => 
                           n5065, ZN => n10163);
   U11359 : NAND3_X1 port map( A1 => n10167, A2 => n10168, A3 => n10169, ZN => 
                           n12076);
   U11360 : AOI221_X1 port map( B1 => n10084, B2 => n5069, C1 => n172, C2 => 
                           MEM_IN(20), A => n10170, ZN => n10169);
   U11361 : OAI22_X1 port map( A1 => n10713, A2 => n273, B1 => n5071, B2 => 
                           n127, ZN => n10170);
   U11362 : AOI22_X1 port map( A1 => n10087, A2 => n5072, B1 => n10088, B2 => 
                           n5073, ZN => n10168);
   U11363 : AOI22_X1 port map( A1 => n10089, A2 => n5074, B1 => n10090, B2 => 
                           n5075, ZN => n10167);
   U11364 : NAND3_X1 port map( A1 => n10171, A2 => n10172, A3 => n10173, ZN => 
                           n12075);
   U11365 : AOI221_X1 port map( B1 => n10084, B2 => n5079, C1 => n172, C2 => 
                           MEM_IN(21), A => n10174, ZN => n10173);
   U11366 : OAI22_X1 port map( A1 => n10712, A2 => n273, B1 => n5081, B2 => 
                           n127, ZN => n10174);
   U11367 : AOI22_X1 port map( A1 => n10087, A2 => n5082, B1 => n10088, B2 => 
                           n5083, ZN => n10172);
   U11368 : AOI22_X1 port map( A1 => n10089, A2 => n5084, B1 => n10090, B2 => 
                           n5085, ZN => n10171);
   U11369 : NAND3_X1 port map( A1 => n10175, A2 => n10176, A3 => n10177, ZN => 
                           n12074);
   U11370 : AOI221_X1 port map( B1 => n10084, B2 => n5089, C1 => n172, C2 => 
                           MEM_IN(22), A => n10178, ZN => n10177);
   U11371 : OAI22_X1 port map( A1 => n10711, A2 => n273, B1 => n5091, B2 => 
                           n127, ZN => n10178);
   U11372 : AOI22_X1 port map( A1 => n10087, A2 => n5092, B1 => n10088, B2 => 
                           n5093, ZN => n10176);
   U11373 : AOI22_X1 port map( A1 => n10089, A2 => n5094, B1 => n10090, B2 => 
                           n5095, ZN => n10175);
   U11374 : NAND3_X1 port map( A1 => n10179, A2 => n10180, A3 => n10181, ZN => 
                           n12073);
   U11375 : AOI221_X1 port map( B1 => n10084, B2 => n5099, C1 => n172, C2 => 
                           MEM_IN(23), A => n10182, ZN => n10181);
   U11376 : OAI22_X1 port map( A1 => n10710, A2 => n273, B1 => n5101, B2 => 
                           n127, ZN => n10182);
   U11377 : AOI22_X1 port map( A1 => n10087, A2 => n5102, B1 => n10088, B2 => 
                           n5103, ZN => n10180);
   U11378 : AOI22_X1 port map( A1 => n10089, A2 => n5104, B1 => n10090, B2 => 
                           n5105, ZN => n10179);
   U11379 : NAND3_X1 port map( A1 => n10183, A2 => n10184, A3 => n10185, ZN => 
                           n12072);
   U11380 : AOI221_X1 port map( B1 => n10084, B2 => n5109, C1 => n172, C2 => 
                           MEM_IN(24), A => n10186, ZN => n10185);
   U11381 : OAI22_X1 port map( A1 => n10709, A2 => n273, B1 => n5111, B2 => 
                           n127, ZN => n10186);
   U11382 : AOI22_X1 port map( A1 => n10087, A2 => n5112, B1 => n10088, B2 => 
                           n5113, ZN => n10184);
   U11383 : AOI22_X1 port map( A1 => n10089, A2 => n5114, B1 => n10090, B2 => 
                           n5115, ZN => n10183);
   U11384 : NAND3_X1 port map( A1 => n10187, A2 => n10188, A3 => n10189, ZN => 
                           n12071);
   U11385 : AOI221_X1 port map( B1 => n10084, B2 => n5119, C1 => n172, C2 => 
                           MEM_IN(25), A => n10190, ZN => n10189);
   U11386 : OAI22_X1 port map( A1 => n10708, A2 => n273, B1 => n5121, B2 => 
                           n127, ZN => n10190);
   U11387 : AOI22_X1 port map( A1 => n10087, A2 => n5122, B1 => n10088, B2 => 
                           n5123, ZN => n10188);
   U11388 : AOI22_X1 port map( A1 => n10089, A2 => n5124, B1 => n10090, B2 => 
                           n5125, ZN => n10187);
   U11389 : NAND3_X1 port map( A1 => n10191, A2 => n10192, A3 => n10193, ZN => 
                           n12070);
   U11390 : AOI221_X1 port map( B1 => n10084, B2 => n5129, C1 => n172, C2 => 
                           MEM_IN(26), A => n10194, ZN => n10193);
   U11391 : OAI22_X1 port map( A1 => n10707, A2 => n273, B1 => n5131, B2 => 
                           n127, ZN => n10194);
   U11392 : AOI22_X1 port map( A1 => n10087, A2 => n5132, B1 => n10088, B2 => 
                           n5133, ZN => n10192);
   U11393 : AOI22_X1 port map( A1 => n10089, A2 => n5134, B1 => n10090, B2 => 
                           n5135, ZN => n10191);
   U11394 : NAND3_X1 port map( A1 => n10195, A2 => n10196, A3 => n10197, ZN => 
                           n12069);
   U11395 : AOI221_X1 port map( B1 => n10084, B2 => n5139, C1 => n172, C2 => 
                           MEM_IN(27), A => n10198, ZN => n10197);
   U11396 : OAI22_X1 port map( A1 => n10706, A2 => n273, B1 => n5141, B2 => 
                           n127, ZN => n10198);
   U11397 : AOI22_X1 port map( A1 => n10087, A2 => n5142, B1 => n10088, B2 => 
                           n5143, ZN => n10196);
   U11398 : AOI22_X1 port map( A1 => n10089, A2 => n5144, B1 => n10090, B2 => 
                           n5145, ZN => n10195);
   U11399 : NAND3_X1 port map( A1 => n10199, A2 => n10200, A3 => n10201, ZN => 
                           n12068);
   U11400 : AOI221_X1 port map( B1 => n10084, B2 => n5149, C1 => n172, C2 => 
                           MEM_IN(28), A => n10202, ZN => n10201);
   U11401 : OAI22_X1 port map( A1 => n10705, A2 => n273, B1 => n5151, B2 => 
                           n127, ZN => n10202);
   U11402 : AOI22_X1 port map( A1 => n10087, A2 => n5152, B1 => n10088, B2 => 
                           n5153, ZN => n10200);
   U11403 : AOI22_X1 port map( A1 => n10089, A2 => n5154, B1 => n10090, B2 => 
                           n5155, ZN => n10199);
   U11404 : NAND3_X1 port map( A1 => n10203, A2 => n10204, A3 => n10205, ZN => 
                           n12067);
   U11405 : AOI221_X1 port map( B1 => n10084, B2 => n5159, C1 => n172, C2 => 
                           MEM_IN(29), A => n10206, ZN => n10205);
   U11406 : OAI22_X1 port map( A1 => n10704, A2 => n273, B1 => n5161, B2 => 
                           n127, ZN => n10206);
   U11407 : AOI22_X1 port map( A1 => n10087, A2 => n5162, B1 => n10088, B2 => 
                           n5163, ZN => n10204);
   U11408 : AOI22_X1 port map( A1 => n10089, A2 => n5164, B1 => n10090, B2 => 
                           n5165, ZN => n10203);
   U11409 : NAND3_X1 port map( A1 => n10207, A2 => n10208, A3 => n10209, ZN => 
                           n12066);
   U11410 : AOI221_X1 port map( B1 => n10084, B2 => n5169, C1 => n172, C2 => 
                           MEM_IN(30), A => n10210, ZN => n10209);
   U11411 : OAI22_X1 port map( A1 => n10703, A2 => n273, B1 => n5171, B2 => 
                           n127, ZN => n10210);
   U11412 : AOI22_X1 port map( A1 => n10087, A2 => n5172, B1 => n10088, B2 => 
                           n5173, ZN => n10208);
   U11413 : AOI22_X1 port map( A1 => n10089, A2 => n5174, B1 => n10090, B2 => 
                           n5175, ZN => n10207);
   U11414 : NAND3_X1 port map( A1 => n10211, A2 => n10212, A3 => n10213, ZN => 
                           n12065);
   U11415 : AOI221_X1 port map( B1 => n10084, B2 => n5179, C1 => n172, C2 => 
                           MEM_IN(31), A => n10214, ZN => n10213);
   U11416 : OAI22_X1 port map( A1 => n10702, A2 => n273, B1 => n5181, B2 => 
                           n127, ZN => n10214);
   U11417 : NAND2_X1 port map( A1 => n5206, A2 => n9921, ZN => n9916);
   U11418 : NAND2_X1 port map( A1 => n9628, A2 => n5206, ZN => n9921);
   U11419 : AOI22_X1 port map( A1 => n10087, A2 => n5191, B1 => n10088, B2 => 
                           n5192, ZN => n10212);
   U11420 : AOI22_X1 port map( A1 => n10089, A2 => n5195, B1 => n10090, B2 => 
                           n5196, ZN => n10211);
   U11421 : OAI22_X1 port map( A1 => n10221, A2 => n10216, B1 => n208, B2 => 
                           n272, ZN => n10218);
   U11422 : NAND3_X1 port map( A1 => n208, A2 => n273, A3 => n9191, ZN => 
                           n10216);
   U11423 : INV_X1 port map( A => n10215, ZN => n9191);
   U11424 : OAI22_X1 port map( A1 => n4786, A2 => n10222, B1 => n10223, B2 => 
                           n5204, ZN => n10086);
   U11425 : NOR2_X1 port map( A1 => n10215, A2 => n10221, ZN => n10223);
   U11426 : NAND2_X1 port map( A1 => n10224, A2 => n9775, ZN => n10215);
   U11427 : AOI211_X1 port map( C1 => n10073, C2 => n5365, A => n10074, B => 
                           n10220, ZN => n10222);
   U11428 : OAI21_X1 port map( B1 => n9775, B2 => n4787, A => n5368, ZN => 
                           n10074);
   U11429 : AND2_X1 port map( A1 => n9628, A2 => n9631, ZN => n9775);
   U11430 : AND2_X1 port map( A1 => n9484, A2 => n9339, ZN => n9628);
   U11431 : NOR3_X1 port map( A1 => n10075, A2 => n10225, A3 => n10076, ZN => 
                           n5365);
   U11432 : INV_X1 port map( A => n10217, ZN => n10221);
   U11433 : AOI21_X1 port map( B1 => n6079, B2 => n10226, A => n10078, ZN => 
                           n10217);
   U11434 : NOR2_X1 port map( A1 => n9339, A2 => n4787, ZN => n9772);
   U11435 : NAND2_X1 port map( A1 => n10080, A2 => n5372, ZN => n9339);
   U11436 : NAND3_X1 port map( A1 => n10227, A2 => n10228, A3 => n10229, ZN => 
                           n12064);
   U11437 : AOI221_X1 port map( B1 => n213, B2 => n4863, C1 => n173, C2 => 
                           MEM_IN(0), A => n10230, ZN => n10229);
   U11438 : OAI22_X1 port map( A1 => n10701, A2 => n259, B1 => n4867, B2 => 
                           n124, ZN => n10230);
   U11439 : AOI22_X1 port map( A1 => n196, A2 => n4869, B1 => n155, B2 => n4871
                           , ZN => n10228);
   U11440 : AOI22_X1 port map( A1 => n239, A2 => n4873, B1 => n152, B2 => n4875
                           , ZN => n10227);
   U11441 : NAND3_X1 port map( A1 => n10232, A2 => n10233, A3 => n10234, ZN => 
                           n12063);
   U11442 : AOI221_X1 port map( B1 => n213, B2 => n4879, C1 => n173, C2 => 
                           MEM_IN(1), A => n10235, ZN => n10234);
   U11443 : OAI22_X1 port map( A1 => n10700, A2 => n259, B1 => n4881, B2 => 
                           n124, ZN => n10235);
   U11444 : AOI22_X1 port map( A1 => n196, A2 => n4882, B1 => n155, B2 => n4883
                           , ZN => n10233);
   U11445 : AOI22_X1 port map( A1 => n239, A2 => n4884, B1 => n152, B2 => n4885
                           , ZN => n10232);
   U11446 : NAND3_X1 port map( A1 => n10236, A2 => n10237, A3 => n10238, ZN => 
                           n12062);
   U11447 : AOI221_X1 port map( B1 => n213, B2 => n4889, C1 => n173, C2 => 
                           MEM_IN(2), A => n10239, ZN => n10238);
   U11448 : OAI22_X1 port map( A1 => n10699, A2 => n259, B1 => n4891, B2 => 
                           n124, ZN => n10239);
   U11449 : AOI22_X1 port map( A1 => n196, A2 => n4892, B1 => n155, B2 => n4893
                           , ZN => n10237);
   U11450 : AOI22_X1 port map( A1 => n239, A2 => n4894, B1 => n152, B2 => n4895
                           , ZN => n10236);
   U11451 : NAND3_X1 port map( A1 => n10240, A2 => n10241, A3 => n10242, ZN => 
                           n12061);
   U11452 : AOI221_X1 port map( B1 => n213, B2 => n4899, C1 => n173, C2 => 
                           MEM_IN(3), A => n10243, ZN => n10242);
   U11453 : OAI22_X1 port map( A1 => n10698, A2 => n259, B1 => n4901, B2 => 
                           n124, ZN => n10243);
   U11454 : AOI22_X1 port map( A1 => n196, A2 => n4902, B1 => n155, B2 => n4903
                           , ZN => n10241);
   U11455 : AOI22_X1 port map( A1 => n239, A2 => n4904, B1 => n152, B2 => n4905
                           , ZN => n10240);
   U11456 : NAND3_X1 port map( A1 => n10244, A2 => n10245, A3 => n10246, ZN => 
                           n12060);
   U11457 : AOI221_X1 port map( B1 => n213, B2 => n4909, C1 => n173, C2 => 
                           MEM_IN(4), A => n10247, ZN => n10246);
   U11458 : OAI22_X1 port map( A1 => n10697, A2 => n259, B1 => n4911, B2 => 
                           n124, ZN => n10247);
   U11459 : AOI22_X1 port map( A1 => n196, A2 => n4912, B1 => n155, B2 => n4913
                           , ZN => n10245);
   U11460 : AOI22_X1 port map( A1 => n239, A2 => n4914, B1 => n152, B2 => n4915
                           , ZN => n10244);
   U11461 : NAND3_X1 port map( A1 => n10248, A2 => n10249, A3 => n10250, ZN => 
                           n12059);
   U11462 : AOI221_X1 port map( B1 => n213, B2 => n4919, C1 => n173, C2 => 
                           MEM_IN(5), A => n10251, ZN => n10250);
   U11463 : OAI22_X1 port map( A1 => n10696, A2 => n259, B1 => n4921, B2 => 
                           n124, ZN => n10251);
   U11464 : AOI22_X1 port map( A1 => n196, A2 => n4922, B1 => n155, B2 => n4923
                           , ZN => n10249);
   U11465 : AOI22_X1 port map( A1 => n239, A2 => n4924, B1 => n152, B2 => n4925
                           , ZN => n10248);
   U11466 : NAND3_X1 port map( A1 => n10252, A2 => n10253, A3 => n10254, ZN => 
                           n12058);
   U11467 : AOI221_X1 port map( B1 => n213, B2 => n4929, C1 => n173, C2 => 
                           MEM_IN(6), A => n10255, ZN => n10254);
   U11468 : OAI22_X1 port map( A1 => n10695, A2 => n259, B1 => n4931, B2 => 
                           n124, ZN => n10255);
   U11469 : AOI22_X1 port map( A1 => n196, A2 => n4932, B1 => n155, B2 => n4933
                           , ZN => n10253);
   U11470 : AOI22_X1 port map( A1 => n239, A2 => n4934, B1 => n152, B2 => n4935
                           , ZN => n10252);
   U11471 : NAND3_X1 port map( A1 => n10256, A2 => n10257, A3 => n10258, ZN => 
                           n12057);
   U11472 : AOI221_X1 port map( B1 => n213, B2 => n4939, C1 => n173, C2 => 
                           MEM_IN(7), A => n10259, ZN => n10258);
   U11473 : OAI22_X1 port map( A1 => n10694, A2 => n259, B1 => n4941, B2 => 
                           n124, ZN => n10259);
   U11474 : AOI22_X1 port map( A1 => n196, A2 => n4942, B1 => n155, B2 => n4943
                           , ZN => n10257);
   U11475 : AOI22_X1 port map( A1 => n239, A2 => n4944, B1 => n152, B2 => n4945
                           , ZN => n10256);
   U11476 : NAND3_X1 port map( A1 => n10260, A2 => n10261, A3 => n10262, ZN => 
                           n12056);
   U11477 : AOI221_X1 port map( B1 => n213, B2 => n4949, C1 => n173, C2 => 
                           MEM_IN(8), A => n10263, ZN => n10262);
   U11478 : OAI22_X1 port map( A1 => n10693, A2 => n259, B1 => n4951, B2 => 
                           n124, ZN => n10263);
   U11479 : AOI22_X1 port map( A1 => n196, A2 => n4952, B1 => n155, B2 => n4953
                           , ZN => n10261);
   U11480 : AOI22_X1 port map( A1 => n239, A2 => n4954, B1 => n152, B2 => n4955
                           , ZN => n10260);
   U11481 : NAND3_X1 port map( A1 => n10264, A2 => n10265, A3 => n10266, ZN => 
                           n12055);
   U11482 : AOI221_X1 port map( B1 => n213, B2 => n4959, C1 => n173, C2 => 
                           MEM_IN(9), A => n10267, ZN => n10266);
   U11483 : OAI22_X1 port map( A1 => n10692, A2 => n259, B1 => n4961, B2 => 
                           n124, ZN => n10267);
   U11484 : AOI22_X1 port map( A1 => n196, A2 => n4962, B1 => n155, B2 => n4963
                           , ZN => n10265);
   U11485 : AOI22_X1 port map( A1 => n239, A2 => n4964, B1 => n152, B2 => n4965
                           , ZN => n10264);
   U11486 : NAND3_X1 port map( A1 => n10268, A2 => n10269, A3 => n10270, ZN => 
                           n12054);
   U11487 : AOI221_X1 port map( B1 => n213, B2 => n4969, C1 => n173, C2 => 
                           MEM_IN(10), A => n10271, ZN => n10270);
   U11488 : OAI22_X1 port map( A1 => n10691, A2 => n259, B1 => n4971, B2 => 
                           n124, ZN => n10271);
   U11489 : AOI22_X1 port map( A1 => n196, A2 => n4972, B1 => n155, B2 => n4973
                           , ZN => n10269);
   U11490 : AOI22_X1 port map( A1 => n239, A2 => n4974, B1 => n152, B2 => n4975
                           , ZN => n10268);
   U11491 : NAND3_X1 port map( A1 => n10272, A2 => n10273, A3 => n10274, ZN => 
                           n12053);
   U11492 : AOI221_X1 port map( B1 => n213, B2 => n4979, C1 => n173, C2 => 
                           MEM_IN(11), A => n10275, ZN => n10274);
   U11493 : OAI22_X1 port map( A1 => n10690, A2 => n259, B1 => n4981, B2 => 
                           n124, ZN => n10275);
   U11494 : AOI22_X1 port map( A1 => n196, A2 => n4982, B1 => n155, B2 => n4983
                           , ZN => n10273);
   U11495 : AOI22_X1 port map( A1 => n239, A2 => n4984, B1 => n152, B2 => n4985
                           , ZN => n10272);
   U11496 : NAND3_X1 port map( A1 => n10276, A2 => n10277, A3 => n10278, ZN => 
                           n12052);
   U11497 : AOI221_X1 port map( B1 => n213, B2 => n4989, C1 => n173, C2 => 
                           MEM_IN(12), A => n10279, ZN => n10278);
   U11498 : OAI22_X1 port map( A1 => n10689, A2 => n259, B1 => n4991, B2 => 
                           n124, ZN => n10279);
   U11499 : AOI22_X1 port map( A1 => n196, A2 => n4992, B1 => n155, B2 => n4993
                           , ZN => n10277);
   U11500 : AOI22_X1 port map( A1 => n239, A2 => n4994, B1 => n152, B2 => n4995
                           , ZN => n10276);
   U11501 : NAND3_X1 port map( A1 => n10280, A2 => n10281, A3 => n10282, ZN => 
                           n12051);
   U11502 : AOI221_X1 port map( B1 => n213, B2 => n4999, C1 => n173, C2 => 
                           MEM_IN(13), A => n10283, ZN => n10282);
   U11503 : OAI22_X1 port map( A1 => n10688, A2 => n259, B1 => n5001, B2 => 
                           n124, ZN => n10283);
   U11504 : AOI22_X1 port map( A1 => n196, A2 => n5002, B1 => n155, B2 => n5003
                           , ZN => n10281);
   U11505 : AOI22_X1 port map( A1 => n239, A2 => n5004, B1 => n152, B2 => n5005
                           , ZN => n10280);
   U11506 : NAND3_X1 port map( A1 => n10284, A2 => n10285, A3 => n10286, ZN => 
                           n12050);
   U11507 : AOI221_X1 port map( B1 => n213, B2 => n5009, C1 => n173, C2 => 
                           MEM_IN(14), A => n10287, ZN => n10286);
   U11508 : OAI22_X1 port map( A1 => n10687, A2 => n259, B1 => n5011, B2 => 
                           n124, ZN => n10287);
   U11509 : AOI22_X1 port map( A1 => n196, A2 => n5012, B1 => n155, B2 => n5013
                           , ZN => n10285);
   U11510 : AOI22_X1 port map( A1 => n239, A2 => n5014, B1 => n152, B2 => n5015
                           , ZN => n10284);
   U11511 : NAND3_X1 port map( A1 => n10288, A2 => n10289, A3 => n10290, ZN => 
                           n12049);
   U11512 : AOI221_X1 port map( B1 => n213, B2 => n5019, C1 => n173, C2 => 
                           MEM_IN(15), A => n10291, ZN => n10290);
   U11513 : OAI22_X1 port map( A1 => n10686, A2 => n259, B1 => n5021, B2 => 
                           n124, ZN => n10291);
   U11514 : AOI22_X1 port map( A1 => n196, A2 => n5022, B1 => n155, B2 => n5023
                           , ZN => n10289);
   U11515 : AOI22_X1 port map( A1 => n239, A2 => n5024, B1 => n152, B2 => n5025
                           , ZN => n10288);
   U11516 : NAND3_X1 port map( A1 => n10292, A2 => n10293, A3 => n10294, ZN => 
                           n12048);
   U11517 : AOI221_X1 port map( B1 => n213, B2 => n5029, C1 => n173, C2 => 
                           MEM_IN(16), A => n10295, ZN => n10294);
   U11518 : OAI22_X1 port map( A1 => n10685, A2 => n259, B1 => n5031, B2 => 
                           n124, ZN => n10295);
   U11519 : AOI22_X1 port map( A1 => n196, A2 => n5032, B1 => n155, B2 => n5033
                           , ZN => n10293);
   U11520 : AOI22_X1 port map( A1 => n239, A2 => n5034, B1 => n152, B2 => n5035
                           , ZN => n10292);
   U11521 : NAND3_X1 port map( A1 => n10296, A2 => n10297, A3 => n10298, ZN => 
                           n12047);
   U11522 : AOI221_X1 port map( B1 => n213, B2 => n5039, C1 => n173, C2 => 
                           MEM_IN(17), A => n10299, ZN => n10298);
   U11523 : OAI22_X1 port map( A1 => n10684, A2 => n259, B1 => n5041, B2 => 
                           n124, ZN => n10299);
   U11524 : AOI22_X1 port map( A1 => n196, A2 => n5042, B1 => n155, B2 => n5043
                           , ZN => n10297);
   U11525 : AOI22_X1 port map( A1 => n239, A2 => n5044, B1 => n152, B2 => n5045
                           , ZN => n10296);
   U11526 : NAND3_X1 port map( A1 => n10300, A2 => n10301, A3 => n10302, ZN => 
                           n12046);
   U11527 : AOI221_X1 port map( B1 => n213, B2 => n5049, C1 => n173, C2 => 
                           MEM_IN(18), A => n10303, ZN => n10302);
   U11528 : OAI22_X1 port map( A1 => n10683, A2 => n259, B1 => n5051, B2 => 
                           n124, ZN => n10303);
   U11529 : AOI22_X1 port map( A1 => n196, A2 => n5052, B1 => n155, B2 => n5053
                           , ZN => n10301);
   U11530 : AOI22_X1 port map( A1 => n239, A2 => n5054, B1 => n152, B2 => n5055
                           , ZN => n10300);
   U11531 : NAND3_X1 port map( A1 => n10304, A2 => n10305, A3 => n10306, ZN => 
                           n12045);
   U11532 : AOI221_X1 port map( B1 => n213, B2 => n5059, C1 => n173, C2 => 
                           MEM_IN(19), A => n10307, ZN => n10306);
   U11533 : OAI22_X1 port map( A1 => n10682, A2 => n259, B1 => n5061, B2 => 
                           n124, ZN => n10307);
   U11534 : AOI22_X1 port map( A1 => n196, A2 => n5062, B1 => n155, B2 => n5063
                           , ZN => n10305);
   U11535 : AOI22_X1 port map( A1 => n239, A2 => n5064, B1 => n152, B2 => n5065
                           , ZN => n10304);
   U11536 : NAND3_X1 port map( A1 => n10308, A2 => n10309, A3 => n10310, ZN => 
                           n12044);
   U11537 : AOI221_X1 port map( B1 => n213, B2 => n5069, C1 => n173, C2 => 
                           MEM_IN(20), A => n10311, ZN => n10310);
   U11538 : OAI22_X1 port map( A1 => n10681, A2 => n259, B1 => n5071, B2 => 
                           n124, ZN => n10311);
   U11539 : AOI22_X1 port map( A1 => n196, A2 => n5072, B1 => n155, B2 => n5073
                           , ZN => n10309);
   U11540 : AOI22_X1 port map( A1 => n239, A2 => n5074, B1 => n152, B2 => n5075
                           , ZN => n10308);
   U11541 : NAND3_X1 port map( A1 => n10312, A2 => n10313, A3 => n10314, ZN => 
                           n12043);
   U11542 : AOI221_X1 port map( B1 => n213, B2 => n5079, C1 => n173, C2 => 
                           MEM_IN(21), A => n10315, ZN => n10314);
   U11543 : OAI22_X1 port map( A1 => n10680, A2 => n259, B1 => n5081, B2 => 
                           n124, ZN => n10315);
   U11544 : AOI22_X1 port map( A1 => n196, A2 => n5082, B1 => n155, B2 => n5083
                           , ZN => n10313);
   U11545 : AOI22_X1 port map( A1 => n239, A2 => n5084, B1 => n152, B2 => n5085
                           , ZN => n10312);
   U11546 : NAND3_X1 port map( A1 => n10316, A2 => n10317, A3 => n10318, ZN => 
                           n12042);
   U11547 : AOI221_X1 port map( B1 => n213, B2 => n5089, C1 => n173, C2 => 
                           MEM_IN(22), A => n10319, ZN => n10318);
   U11548 : OAI22_X1 port map( A1 => n10679, A2 => n259, B1 => n5091, B2 => 
                           n124, ZN => n10319);
   U11549 : AOI22_X1 port map( A1 => n196, A2 => n5092, B1 => n155, B2 => n5093
                           , ZN => n10317);
   U11550 : AOI22_X1 port map( A1 => n239, A2 => n5094, B1 => n152, B2 => n5095
                           , ZN => n10316);
   U11551 : NAND3_X1 port map( A1 => n10320, A2 => n10321, A3 => n10322, ZN => 
                           n12041);
   U11552 : AOI221_X1 port map( B1 => n213, B2 => n5099, C1 => n173, C2 => 
                           MEM_IN(23), A => n10387, ZN => n10322);
   U11553 : OAI22_X1 port map( A1 => n10678, A2 => n259, B1 => n5101, B2 => 
                           n124, ZN => n10387);
   U11554 : AOI22_X1 port map( A1 => n196, A2 => n5102, B1 => n155, B2 => n5103
                           , ZN => n10321);
   U11555 : AOI22_X1 port map( A1 => n239, A2 => n5104, B1 => n152, B2 => n5105
                           , ZN => n10320);
   U11556 : NAND3_X1 port map( A1 => n10414, A2 => n10415, A3 => n10416, ZN => 
                           n12040);
   U11557 : AOI221_X1 port map( B1 => n213, B2 => n5109, C1 => n173, C2 => 
                           MEM_IN(24), A => n10417, ZN => n10416);
   U11558 : OAI22_X1 port map( A1 => n10677, A2 => n259, B1 => n5111, B2 => 
                           n124, ZN => n10417);
   U11559 : AOI22_X1 port map( A1 => n196, A2 => n5112, B1 => n155, B2 => n5113
                           , ZN => n10415);
   U11560 : AOI22_X1 port map( A1 => n239, A2 => n5114, B1 => n152, B2 => n5115
                           , ZN => n10414);
   U11561 : NAND3_X1 port map( A1 => n10418, A2 => n10419, A3 => n10420, ZN => 
                           n12039);
   U11562 : AOI221_X1 port map( B1 => n213, B2 => n5119, C1 => n173, C2 => 
                           MEM_IN(25), A => n10421, ZN => n10420);
   U11563 : OAI22_X1 port map( A1 => n10676, A2 => n259, B1 => n5121, B2 => 
                           n124, ZN => n10421);
   U11564 : AOI22_X1 port map( A1 => n196, A2 => n5122, B1 => n155, B2 => n5123
                           , ZN => n10419);
   U11565 : AOI22_X1 port map( A1 => n239, A2 => n5124, B1 => n152, B2 => n5125
                           , ZN => n10418);
   U11566 : NAND3_X1 port map( A1 => n10422, A2 => n10423, A3 => n10424, ZN => 
                           n12038);
   U11567 : AOI221_X1 port map( B1 => n213, B2 => n5129, C1 => n173, C2 => 
                           MEM_IN(26), A => n10425, ZN => n10424);
   U11568 : OAI22_X1 port map( A1 => n10675, A2 => n259, B1 => n5131, B2 => 
                           n124, ZN => n10425);
   U11569 : AOI22_X1 port map( A1 => n196, A2 => n5132, B1 => n155, B2 => n5133
                           , ZN => n10423);
   U11570 : AOI22_X1 port map( A1 => n239, A2 => n5134, B1 => n152, B2 => n5135
                           , ZN => n10422);
   U11571 : NAND3_X1 port map( A1 => n10426, A2 => n10427, A3 => n10428, ZN => 
                           n12037);
   U11572 : AOI221_X1 port map( B1 => n213, B2 => n5139, C1 => n173, C2 => 
                           MEM_IN(27), A => n10429, ZN => n10428);
   U11573 : OAI22_X1 port map( A1 => n10674, A2 => n259, B1 => n5141, B2 => 
                           n124, ZN => n10429);
   U11574 : AOI22_X1 port map( A1 => n196, A2 => n5142, B1 => n155, B2 => n5143
                           , ZN => n10427);
   U11575 : AOI22_X1 port map( A1 => n239, A2 => n5144, B1 => n152, B2 => n5145
                           , ZN => n10426);
   U11576 : NAND3_X1 port map( A1 => n10430, A2 => n10431, A3 => n10432, ZN => 
                           n12036);
   U11577 : AOI221_X1 port map( B1 => n213, B2 => n5149, C1 => n173, C2 => 
                           MEM_IN(28), A => n10433, ZN => n10432);
   U11578 : OAI22_X1 port map( A1 => n10673, A2 => n259, B1 => n5151, B2 => 
                           n124, ZN => n10433);
   U11579 : AOI22_X1 port map( A1 => n196, A2 => n5152, B1 => n155, B2 => n5153
                           , ZN => n10431);
   U11580 : AOI22_X1 port map( A1 => n239, A2 => n5154, B1 => n152, B2 => n5155
                           , ZN => n10430);
   U11581 : NAND3_X1 port map( A1 => n10434, A2 => n10435, A3 => n10436, ZN => 
                           n12035);
   U11582 : AOI221_X1 port map( B1 => n213, B2 => n5159, C1 => n173, C2 => 
                           MEM_IN(29), A => n10437, ZN => n10436);
   U11583 : OAI22_X1 port map( A1 => n10672, A2 => n259, B1 => n5161, B2 => 
                           n124, ZN => n10437);
   U11584 : AOI22_X1 port map( A1 => n196, A2 => n5162, B1 => n155, B2 => n5163
                           , ZN => n10435);
   U11585 : AOI22_X1 port map( A1 => n239, A2 => n5164, B1 => n152, B2 => n5165
                           , ZN => n10434);
   U11586 : NAND3_X1 port map( A1 => n10438, A2 => n10439, A3 => n10440, ZN => 
                           n12034);
   U11587 : AOI221_X1 port map( B1 => n213, B2 => n5169, C1 => n173, C2 => 
                           MEM_IN(30), A => n10441, ZN => n10440);
   U11588 : OAI22_X1 port map( A1 => n10671, A2 => n259, B1 => n5171, B2 => 
                           n124, ZN => n10441);
   U11589 : AOI22_X1 port map( A1 => n196, A2 => n5172, B1 => n155, B2 => n5173
                           , ZN => n10439);
   U11590 : AOI22_X1 port map( A1 => n239, A2 => n5174, B1 => n152, B2 => n5175
                           , ZN => n10438);
   U11591 : NAND3_X1 port map( A1 => n10442, A2 => n10443, A3 => n10444, ZN => 
                           n12033);
   U11592 : AOI221_X1 port map( B1 => n213, B2 => n5179, C1 => n173, C2 => 
                           MEM_IN(31), A => n10445, ZN => n10444);
   U11593 : OAI22_X1 port map( A1 => n10670, A2 => n259, B1 => n5181, B2 => 
                           n124, ZN => n10445);
   U11594 : INV_X1 port map( A => n11848, ZN => n11847);
   U11595 : AOI22_X1 port map( A1 => n196, A2 => n5191, B1 => n155, B2 => n5192
                           , ZN => n10443);
   U11596 : AOI22_X1 port map( A1 => n239, A2 => n5195, B1 => n152, B2 => n5196
                           , ZN => n10442);
   U11597 : INV_X1 port map( A => n10068, ZN => n10067);
   U11598 : AOI22_X1 port map( A1 => n11845, A2 => n11851, B1 => n4841, B2 => 
                           n259, ZN => n11846);
   U11599 : INV_X1 port map( A => n11844, ZN => n11851);
   U11600 : NAND3_X1 port map( A1 => n208, A2 => n259, A3 => n9338, ZN => 
                           n11844);
   U11601 : INV_X1 port map( A => n11843, ZN => n9338);
   U11602 : OAI22_X1 port map( A1 => n4786, A2 => n11852, B1 => n11853, B2 => 
                           n5204, ZN => n10231);
   U11603 : NOR2_X1 port map( A1 => n11843, A2 => n11854, ZN => n11853);
   U11604 : NAND4_X1 port map( A1 => n10224, A2 => n9631, A3 => n9484, A4 => 
                           n11855, ZN => n11843);
   U11605 : AND4_X1 port map( A1 => n11856, A2 => n10219, A3 => n5368, A4 => 
                           n11849, ZN => n11852);
   U11606 : INV_X1 port map( A => n10220, ZN => n10219);
   U11607 : AOI211_X1 port map( C1 => n5522, C2 => n10073, A => n9918, B => 
                           n10068, ZN => n11856);
   U11608 : NOR2_X1 port map( A1 => n9484, A2 => n4787, ZN => n9918);
   U11609 : NOR3_X1 port map( A1 => n10076, A2 => n11857, A3 => n10077, ZN => 
                           n5522);
   U11610 : INV_X1 port map( A => n11854, ZN => n11845);
   U11611 : NAND3_X1 port map( A1 => n11858, A2 => n11870, A3 => n11871, ZN => 
                           n11854);
   U11612 : NAND2_X1 port map( A1 => n10080, A2 => n5526, ZN => n9484);
   U11613 : NAND3_X1 port map( A1 => n13193, A2 => n13194, A3 => n13195, ZN => 
                           n12032);
   U11614 : AOI221_X1 port map( B1 => n13196, B2 => n4863, C1 => n170, C2 => 
                           MEM_IN(0), A => n13197, ZN => n13195);
   U11615 : OAI22_X1 port map( A1 => n10669, A2 => n275, B1 => n4867, B2 => 
                           n125, ZN => n13197);
   U11616 : AOI22_X1 port map( A1 => n13199, A2 => n4869, B1 => n13200, B2 => 
                           n4871, ZN => n13194);
   U11617 : AOI22_X1 port map( A1 => n13201, A2 => n4873, B1 => n13202, B2 => 
                           n4875, ZN => n13193);
   U11618 : NAND3_X1 port map( A1 => n13203, A2 => n13204, A3 => n13205, ZN => 
                           n12031);
   U11619 : AOI221_X1 port map( B1 => n13196, B2 => n4879, C1 => n170, C2 => 
                           MEM_IN(1), A => n13206, ZN => n13205);
   U11620 : OAI22_X1 port map( A1 => n10668, A2 => n275, B1 => n4881, B2 => 
                           n125, ZN => n13206);
   U11621 : AOI22_X1 port map( A1 => n13199, A2 => n4882, B1 => n13200, B2 => 
                           n4883, ZN => n13204);
   U11622 : AOI22_X1 port map( A1 => n13201, A2 => n4884, B1 => n13202, B2 => 
                           n4885, ZN => n13203);
   U11623 : NAND3_X1 port map( A1 => n13207, A2 => n13208, A3 => n13209, ZN => 
                           n12030);
   U11624 : AOI221_X1 port map( B1 => n13196, B2 => n4889, C1 => n170, C2 => 
                           MEM_IN(2), A => n13210, ZN => n13209);
   U11625 : OAI22_X1 port map( A1 => n10667, A2 => n275, B1 => n4891, B2 => 
                           n125, ZN => n13210);
   U11626 : AOI22_X1 port map( A1 => n13199, A2 => n4892, B1 => n13200, B2 => 
                           n4893, ZN => n13208);
   U11627 : AOI22_X1 port map( A1 => n13201, A2 => n4894, B1 => n13202, B2 => 
                           n4895, ZN => n13207);
   U11628 : NAND3_X1 port map( A1 => n13211, A2 => n13212, A3 => n13213, ZN => 
                           n12029);
   U11629 : AOI221_X1 port map( B1 => n13196, B2 => n4899, C1 => n170, C2 => 
                           MEM_IN(3), A => n13214, ZN => n13213);
   U11630 : OAI22_X1 port map( A1 => n10666, A2 => n275, B1 => n4901, B2 => 
                           n125, ZN => n13214);
   U11631 : AOI22_X1 port map( A1 => n13199, A2 => n4902, B1 => n13200, B2 => 
                           n4903, ZN => n13212);
   U11632 : AOI22_X1 port map( A1 => n13201, A2 => n4904, B1 => n13202, B2 => 
                           n4905, ZN => n13211);
   U11633 : NAND3_X1 port map( A1 => n13215, A2 => n13216, A3 => n13217, ZN => 
                           n12028);
   U11634 : AOI221_X1 port map( B1 => n13196, B2 => n4909, C1 => n170, C2 => 
                           MEM_IN(4), A => n13218, ZN => n13217);
   U11635 : OAI22_X1 port map( A1 => n10665, A2 => n275, B1 => n4911, B2 => 
                           n125, ZN => n13218);
   U11636 : AOI22_X1 port map( A1 => n13199, A2 => n4912, B1 => n13200, B2 => 
                           n4913, ZN => n13216);
   U11637 : AOI22_X1 port map( A1 => n13201, A2 => n4914, B1 => n13202, B2 => 
                           n4915, ZN => n13215);
   U11638 : NAND3_X1 port map( A1 => n13219, A2 => n13220, A3 => n13221, ZN => 
                           n12027);
   U11639 : AOI221_X1 port map( B1 => n13196, B2 => n4919, C1 => n170, C2 => 
                           MEM_IN(5), A => n13222, ZN => n13221);
   U11640 : OAI22_X1 port map( A1 => n10664, A2 => n275, B1 => n4921, B2 => 
                           n125, ZN => n13222);
   U11641 : AOI22_X1 port map( A1 => n13199, A2 => n4922, B1 => n13200, B2 => 
                           n4923, ZN => n13220);
   U11642 : AOI22_X1 port map( A1 => n13201, A2 => n4924, B1 => n13202, B2 => 
                           n4925, ZN => n13219);
   U11643 : NAND3_X1 port map( A1 => n13223, A2 => n13224, A3 => n13225, ZN => 
                           n12026);
   U11644 : AOI221_X1 port map( B1 => n13196, B2 => n4929, C1 => n170, C2 => 
                           MEM_IN(6), A => n13226, ZN => n13225);
   U11645 : OAI22_X1 port map( A1 => n10663, A2 => n275, B1 => n4931, B2 => 
                           n125, ZN => n13226);
   U11646 : AOI22_X1 port map( A1 => n13199, A2 => n4932, B1 => n13200, B2 => 
                           n4933, ZN => n13224);
   U11647 : AOI22_X1 port map( A1 => n13201, A2 => n4934, B1 => n13202, B2 => 
                           n4935, ZN => n13223);
   U11648 : NAND3_X1 port map( A1 => n13227, A2 => n13228, A3 => n13229, ZN => 
                           n12025);
   U11649 : AOI221_X1 port map( B1 => n13196, B2 => n4939, C1 => n170, C2 => 
                           MEM_IN(7), A => n13230, ZN => n13229);
   U11650 : OAI22_X1 port map( A1 => n10662, A2 => n275, B1 => n4941, B2 => 
                           n125, ZN => n13230);
   U11651 : AOI22_X1 port map( A1 => n13199, A2 => n4942, B1 => n13200, B2 => 
                           n4943, ZN => n13228);
   U11652 : AOI22_X1 port map( A1 => n13201, A2 => n4944, B1 => n13202, B2 => 
                           n4945, ZN => n13227);
   U11653 : NAND3_X1 port map( A1 => n13231, A2 => n13232, A3 => n13233, ZN => 
                           n12024);
   U11654 : AOI221_X1 port map( B1 => n13196, B2 => n4949, C1 => n170, C2 => 
                           MEM_IN(8), A => n13234, ZN => n13233);
   U11655 : OAI22_X1 port map( A1 => n10661, A2 => n275, B1 => n4951, B2 => 
                           n125, ZN => n13234);
   U11656 : AOI22_X1 port map( A1 => n13199, A2 => n4952, B1 => n13200, B2 => 
                           n4953, ZN => n13232);
   U11657 : AOI22_X1 port map( A1 => n13201, A2 => n4954, B1 => n13202, B2 => 
                           n4955, ZN => n13231);
   U11658 : NAND3_X1 port map( A1 => n13235, A2 => n13236, A3 => n13237, ZN => 
                           n12023);
   U11659 : AOI221_X1 port map( B1 => n13196, B2 => n4959, C1 => n170, C2 => 
                           MEM_IN(9), A => n13238, ZN => n13237);
   U11660 : OAI22_X1 port map( A1 => n10660, A2 => n275, B1 => n4961, B2 => 
                           n125, ZN => n13238);
   U11661 : AOI22_X1 port map( A1 => n13199, A2 => n4962, B1 => n13200, B2 => 
                           n4963, ZN => n13236);
   U11662 : AOI22_X1 port map( A1 => n13201, A2 => n4964, B1 => n13202, B2 => 
                           n4965, ZN => n13235);
   U11663 : NAND3_X1 port map( A1 => n13239, A2 => n13240, A3 => n13241, ZN => 
                           n12022);
   U11664 : AOI221_X1 port map( B1 => n13196, B2 => n4969, C1 => n170, C2 => 
                           MEM_IN(10), A => n13242, ZN => n13241);
   U11665 : OAI22_X1 port map( A1 => n10659, A2 => n275, B1 => n4971, B2 => 
                           n125, ZN => n13242);
   U11666 : AOI22_X1 port map( A1 => n13199, A2 => n4972, B1 => n13200, B2 => 
                           n4973, ZN => n13240);
   U11667 : AOI22_X1 port map( A1 => n13201, A2 => n4974, B1 => n13202, B2 => 
                           n4975, ZN => n13239);
   U11668 : NAND3_X1 port map( A1 => n13243, A2 => n13244, A3 => n13245, ZN => 
                           n12021);
   U11669 : AOI221_X1 port map( B1 => n13196, B2 => n4979, C1 => n170, C2 => 
                           MEM_IN(11), A => n13246, ZN => n13245);
   U11670 : OAI22_X1 port map( A1 => n10658, A2 => n275, B1 => n4981, B2 => 
                           n125, ZN => n13246);
   U11671 : AOI22_X1 port map( A1 => n13199, A2 => n4982, B1 => n13200, B2 => 
                           n4983, ZN => n13244);
   U11672 : AOI22_X1 port map( A1 => n13201, A2 => n4984, B1 => n13202, B2 => 
                           n4985, ZN => n13243);
   U11673 : NAND3_X1 port map( A1 => n13247, A2 => n13248, A3 => n13249, ZN => 
                           n12020);
   U11674 : AOI221_X1 port map( B1 => n13196, B2 => n4989, C1 => n170, C2 => 
                           MEM_IN(12), A => n13250, ZN => n13249);
   U11675 : OAI22_X1 port map( A1 => n10657, A2 => n275, B1 => n4991, B2 => 
                           n125, ZN => n13250);
   U11676 : AOI22_X1 port map( A1 => n13199, A2 => n4992, B1 => n13200, B2 => 
                           n4993, ZN => n13248);
   U11677 : AOI22_X1 port map( A1 => n13201, A2 => n4994, B1 => n13202, B2 => 
                           n4995, ZN => n13247);
   U11678 : NAND3_X1 port map( A1 => n13251, A2 => n13252, A3 => n13253, ZN => 
                           n12019);
   U11679 : AOI221_X1 port map( B1 => n13196, B2 => n4999, C1 => n170, C2 => 
                           MEM_IN(13), A => n13254, ZN => n13253);
   U11680 : OAI22_X1 port map( A1 => n10656, A2 => n275, B1 => n5001, B2 => 
                           n125, ZN => n13254);
   U11681 : AOI22_X1 port map( A1 => n13199, A2 => n5002, B1 => n13200, B2 => 
                           n5003, ZN => n13252);
   U11682 : AOI22_X1 port map( A1 => n13201, A2 => n5004, B1 => n13202, B2 => 
                           n5005, ZN => n13251);
   U11683 : NAND3_X1 port map( A1 => n13255, A2 => n13256, A3 => n13257, ZN => 
                           n12018);
   U11684 : AOI221_X1 port map( B1 => n13196, B2 => n5009, C1 => n170, C2 => 
                           MEM_IN(14), A => n13258, ZN => n13257);
   U11685 : OAI22_X1 port map( A1 => n10655, A2 => n275, B1 => n5011, B2 => 
                           n125, ZN => n13258);
   U11686 : AOI22_X1 port map( A1 => n13199, A2 => n5012, B1 => n13200, B2 => 
                           n5013, ZN => n13256);
   U11687 : AOI22_X1 port map( A1 => n13201, A2 => n5014, B1 => n13202, B2 => 
                           n5015, ZN => n13255);
   U11688 : NAND3_X1 port map( A1 => n13259, A2 => n13260, A3 => n13261, ZN => 
                           n12017);
   U11689 : AOI221_X1 port map( B1 => n13196, B2 => n5019, C1 => n170, C2 => 
                           MEM_IN(15), A => n13262, ZN => n13261);
   U11690 : OAI22_X1 port map( A1 => n10654, A2 => n275, B1 => n5021, B2 => 
                           n125, ZN => n13262);
   U11691 : AOI22_X1 port map( A1 => n13199, A2 => n5022, B1 => n13200, B2 => 
                           n5023, ZN => n13260);
   U11692 : AOI22_X1 port map( A1 => n13201, A2 => n5024, B1 => n13202, B2 => 
                           n5025, ZN => n13259);
   U11693 : NAND3_X1 port map( A1 => n13263, A2 => n13264, A3 => n13265, ZN => 
                           n12016);
   U11694 : AOI221_X1 port map( B1 => n13196, B2 => n5029, C1 => n170, C2 => 
                           MEM_IN(16), A => n13266, ZN => n13265);
   U11695 : OAI22_X1 port map( A1 => n10653, A2 => n275, B1 => n5031, B2 => 
                           n125, ZN => n13266);
   U11696 : AOI22_X1 port map( A1 => n13199, A2 => n5032, B1 => n13200, B2 => 
                           n5033, ZN => n13264);
   U11697 : AOI22_X1 port map( A1 => n13201, A2 => n5034, B1 => n13202, B2 => 
                           n5035, ZN => n13263);
   U11698 : NAND3_X1 port map( A1 => n13267, A2 => n13268, A3 => n13269, ZN => 
                           n12015);
   U11699 : AOI221_X1 port map( B1 => n13196, B2 => n5039, C1 => n170, C2 => 
                           MEM_IN(17), A => n13270, ZN => n13269);
   U11700 : OAI22_X1 port map( A1 => n10652, A2 => n275, B1 => n5041, B2 => 
                           n125, ZN => n13270);
   U11701 : AOI22_X1 port map( A1 => n13199, A2 => n5042, B1 => n13200, B2 => 
                           n5043, ZN => n13268);
   U11702 : AOI22_X1 port map( A1 => n13201, A2 => n5044, B1 => n13202, B2 => 
                           n5045, ZN => n13267);
   U11703 : NAND3_X1 port map( A1 => n13271, A2 => n13272, A3 => n13273, ZN => 
                           n12014);
   U11704 : AOI221_X1 port map( B1 => n13196, B2 => n5049, C1 => n170, C2 => 
                           MEM_IN(18), A => n13274, ZN => n13273);
   U11705 : OAI22_X1 port map( A1 => n10651, A2 => n275, B1 => n5051, B2 => 
                           n125, ZN => n13274);
   U11706 : AOI22_X1 port map( A1 => n13199, A2 => n5052, B1 => n13200, B2 => 
                           n5053, ZN => n13272);
   U11707 : AOI22_X1 port map( A1 => n13201, A2 => n5054, B1 => n13202, B2 => 
                           n5055, ZN => n13271);
   U11708 : NAND3_X1 port map( A1 => n13275, A2 => n13276, A3 => n13277, ZN => 
                           n12013);
   U11709 : AOI221_X1 port map( B1 => n13196, B2 => n5059, C1 => n170, C2 => 
                           MEM_IN(19), A => n13278, ZN => n13277);
   U11710 : OAI22_X1 port map( A1 => n10650, A2 => n275, B1 => n5061, B2 => 
                           n125, ZN => n13278);
   U11711 : AOI22_X1 port map( A1 => n13199, A2 => n5062, B1 => n13200, B2 => 
                           n5063, ZN => n13276);
   U11712 : AOI22_X1 port map( A1 => n13201, A2 => n5064, B1 => n13202, B2 => 
                           n5065, ZN => n13275);
   U11713 : NAND3_X1 port map( A1 => n13279, A2 => n13280, A3 => n13281, ZN => 
                           n12012);
   U11714 : AOI221_X1 port map( B1 => n13196, B2 => n5069, C1 => n170, C2 => 
                           MEM_IN(20), A => n13282, ZN => n13281);
   U11715 : OAI22_X1 port map( A1 => n10649, A2 => n275, B1 => n5071, B2 => 
                           n125, ZN => n13282);
   U11718 : AOI22_X1 port map( A1 => n13199, A2 => n5072, B1 => n13200, B2 => 
                           n5073, ZN => n13280);
   U11719 : AOI22_X1 port map( A1 => n13201, A2 => n5074, B1 => n13202, B2 => 
                           n5075, ZN => n13279);
   U11721 : NAND3_X1 port map( A1 => n13283, A2 => n13284, A3 => n13285, ZN => 
                           n12011);
   U11722 : AOI221_X1 port map( B1 => n13196, B2 => n5079, C1 => n170, C2 => 
                           MEM_IN(21), A => n13286, ZN => n13285);
   U11723 : OAI22_X1 port map( A1 => n10648, A2 => n275, B1 => n5081, B2 => 
                           n125, ZN => n13286);
   U11724 : AOI22_X1 port map( A1 => n13199, A2 => n5082, B1 => n13200, B2 => 
                           n5083, ZN => n13284);
   U11725 : AOI22_X1 port map( A1 => n13201, A2 => n5084, B1 => n13202, B2 => 
                           n5085, ZN => n13283);
   U11726 : NAND3_X1 port map( A1 => n13287, A2 => n13288, A3 => n13289, ZN => 
                           n12010);
   U11727 : AOI221_X1 port map( B1 => n13196, B2 => n5089, C1 => n170, C2 => 
                           MEM_IN(22), A => n13290, ZN => n13289);
   U11728 : OAI22_X1 port map( A1 => n10647, A2 => n275, B1 => n5091, B2 => 
                           n125, ZN => n13290);
   U11729 : AOI22_X1 port map( A1 => n13199, A2 => n5092, B1 => n13200, B2 => 
                           n5093, ZN => n13288);
   U11730 : AOI22_X1 port map( A1 => n13201, A2 => n5094, B1 => n13202, B2 => 
                           n5095, ZN => n13287);
   U11731 : NAND3_X1 port map( A1 => n13291, A2 => n13292, A3 => n13293, ZN => 
                           n12009);
   U11732 : AOI221_X1 port map( B1 => n13196, B2 => n5099, C1 => n170, C2 => 
                           MEM_IN(23), A => n13294, ZN => n13293);
   U11733 : OAI22_X1 port map( A1 => n10646, A2 => n275, B1 => n5101, B2 => 
                           n125, ZN => n13294);
   U11734 : AOI22_X1 port map( A1 => n13199, A2 => n5102, B1 => n13200, B2 => 
                           n5103, ZN => n13292);
   U11735 : AOI22_X1 port map( A1 => n13201, A2 => n5104, B1 => n13202, B2 => 
                           n5105, ZN => n13291);
   U11736 : NAND3_X1 port map( A1 => n13295, A2 => n13296, A3 => n13297, ZN => 
                           n12008);
   U11737 : AOI221_X1 port map( B1 => n13196, B2 => n5109, C1 => n170, C2 => 
                           MEM_IN(24), A => n13298, ZN => n13297);
   U11738 : OAI22_X1 port map( A1 => n10645, A2 => n275, B1 => n5111, B2 => 
                           n125, ZN => n13298);
   U11739 : AOI22_X1 port map( A1 => n13199, A2 => n5112, B1 => n13200, B2 => 
                           n5113, ZN => n13296);
   U11740 : AOI22_X1 port map( A1 => n13201, A2 => n5114, B1 => n13202, B2 => 
                           n5115, ZN => n13295);
   U11741 : NAND3_X1 port map( A1 => n13299, A2 => n13300, A3 => n13301, ZN => 
                           n12007);
   U11742 : AOI221_X1 port map( B1 => n13196, B2 => n5119, C1 => n170, C2 => 
                           MEM_IN(25), A => n13302, ZN => n13301);
   U11743 : OAI22_X1 port map( A1 => n10644, A2 => n275, B1 => n5121, B2 => 
                           n125, ZN => n13302);
   U11744 : AOI22_X1 port map( A1 => n13199, A2 => n5122, B1 => n13200, B2 => 
                           n5123, ZN => n13300);
   U11745 : AOI22_X1 port map( A1 => n13201, A2 => n5124, B1 => n13202, B2 => 
                           n5125, ZN => n13299);
   U11746 : NAND3_X1 port map( A1 => n13303, A2 => n13304, A3 => n13305, ZN => 
                           n12006);
   U11747 : AOI221_X1 port map( B1 => n13196, B2 => n5129, C1 => n170, C2 => 
                           MEM_IN(26), A => n13306, ZN => n13305);
   U11748 : OAI22_X1 port map( A1 => n10643, A2 => n275, B1 => n5131, B2 => 
                           n125, ZN => n13306);
   U11749 : AOI22_X1 port map( A1 => n13199, A2 => n5132, B1 => n13200, B2 => 
                           n5133, ZN => n13304);
   U11750 : AOI22_X1 port map( A1 => n13201, A2 => n5134, B1 => n13202, B2 => 
                           n5135, ZN => n13303);
   U11751 : NAND3_X1 port map( A1 => n13307, A2 => n13308, A3 => n13309, ZN => 
                           n12005);
   U11752 : AOI221_X1 port map( B1 => n13196, B2 => n5139, C1 => n170, C2 => 
                           MEM_IN(27), A => n13310, ZN => n13309);
   U11753 : OAI22_X1 port map( A1 => n10642, A2 => n275, B1 => n5141, B2 => 
                           n125, ZN => n13310);
   U11754 : AOI22_X1 port map( A1 => n13199, A2 => n5142, B1 => n13200, B2 => 
                           n5143, ZN => n13308);
   U11755 : AOI22_X1 port map( A1 => n13201, A2 => n5144, B1 => n13202, B2 => 
                           n5145, ZN => n13307);
   U11756 : NAND3_X1 port map( A1 => n13311, A2 => n13312, A3 => n13313, ZN => 
                           n12004);
   U11757 : AOI221_X1 port map( B1 => n13196, B2 => n5149, C1 => n170, C2 => 
                           MEM_IN(28), A => n13314, ZN => n13313);
   U11758 : OAI22_X1 port map( A1 => n10641, A2 => n275, B1 => n5151, B2 => 
                           n125, ZN => n13314);
   U11759 : AOI22_X1 port map( A1 => n13199, A2 => n5152, B1 => n13200, B2 => 
                           n5153, ZN => n13312);
   U11760 : AOI22_X1 port map( A1 => n13201, A2 => n5154, B1 => n13202, B2 => 
                           n5155, ZN => n13311);
   U11761 : NAND3_X1 port map( A1 => n13315, A2 => n13316, A3 => n13317, ZN => 
                           n12003);
   U11762 : AOI221_X1 port map( B1 => n13196, B2 => n5159, C1 => n170, C2 => 
                           MEM_IN(29), A => n13318, ZN => n13317);
   U11763 : OAI22_X1 port map( A1 => n10640, A2 => n275, B1 => n5161, B2 => 
                           n125, ZN => n13318);
   U11764 : AOI22_X1 port map( A1 => n13199, A2 => n5162, B1 => n13200, B2 => 
                           n5163, ZN => n13316);
   U11765 : AOI22_X1 port map( A1 => n13201, A2 => n5164, B1 => n13202, B2 => 
                           n5165, ZN => n13315);
   U11766 : NAND3_X1 port map( A1 => n13319, A2 => n13320, A3 => n13321, ZN => 
                           n12002);
   U11767 : AOI221_X1 port map( B1 => n13196, B2 => n5169, C1 => n170, C2 => 
                           MEM_IN(30), A => n13322, ZN => n13321);
   U11768 : OAI22_X1 port map( A1 => n10639, A2 => n275, B1 => n5171, B2 => 
                           n125, ZN => n13322);
   U11769 : AOI22_X1 port map( A1 => n13199, A2 => n5172, B1 => n13200, B2 => 
                           n5173, ZN => n13320);
   U11770 : AOI22_X1 port map( A1 => n13201, A2 => n5174, B1 => n13202, B2 => 
                           n5175, ZN => n13319);
   U11771 : NAND3_X1 port map( A1 => n13323, A2 => n13324, A3 => n13325, ZN => 
                           n12001);
   U11772 : AOI221_X1 port map( B1 => n13196, B2 => n5179, C1 => n170, C2 => 
                           MEM_IN(31), A => n13326, ZN => n13325);
   U11773 : OAI22_X1 port map( A1 => n10638, A2 => n275, B1 => n5181, B2 => 
                           n125, ZN => n13326);
   U11774 : INV_X1 port map( A => n13330, ZN => n13329);
   U11775 : NAND2_X1 port map( A1 => n5206, A2 => n11850, ZN => n11848);
   U11776 : NAND3_X1 port map( A1 => n5206, A2 => n9631, A3 => n10072, ZN => 
                           n11850);
   U11777 : AOI22_X1 port map( A1 => n13199, A2 => n5191, B1 => n13200, B2 => 
                           n5192, ZN => n13324);
   U11778 : AOI22_X1 port map( A1 => n13201, A2 => n5195, B1 => n13202, B2 => 
                           n5196, ZN => n13323);
   U11779 : OAI22_X1 port map( A1 => n13330, A2 => n13328, B1 => n208, B2 => 
                           n274, ZN => n13332);
   U11780 : NAND3_X1 port map( A1 => n208, A2 => n275, A3 => n9483, ZN => 
                           n13328);
   U11781 : INV_X1 port map( A => n13327, ZN => n9483);
   U11782 : OAI22_X1 port map( A1 => n4786, A2 => n13335, B1 => n13336, B2 => 
                           n5204, ZN => n13198);
   U11783 : NOR2_X1 port map( A1 => n13327, A2 => n13330, ZN => n13336);
   U11784 : NAND3_X1 port map( A1 => n10224, A2 => n9631, A3 => n13337, ZN => 
                           n13327);
   U11785 : NOR3_X1 port map( A1 => n13338, A2 => RESET, A3 => n10068, ZN => 
                           n13335);
   U11786 : OAI22_X1 port map( A1 => n10224, A2 => n4787, B1 => n5771, B2 => 
                           n13339, ZN => n13338);
   U11787 : INV_X1 port map( A => n9337, ZN => n5771);
   U11788 : NOR3_X1 port map( A1 => n11857, A2 => n10225, A3 => n10076, ZN => 
                           n9337);
   U11789 : OAI211_X1 port map( C1 => n13340, C2 => n13341, A => n11870, B => 
                           n11871, ZN => n13330);
   U11790 : INV_X1 port map( A => n6381, ZN => n13340);
   U11791 : NOR2_X1 port map( A1 => n9631, A2 => n4787, ZN => n10068);
   U11792 : NAND2_X1 port map( A1 => n10080, A2 => n5775, ZN => n9631);
   U11793 : NAND3_X1 port map( A1 => n13342, A2 => n13343, A3 => n13344, ZN => 
                           n12000);
   U11794 : AOI221_X1 port map( B1 => n13345, B2 => n4863, C1 => n171, C2 => 
                           MEM_IN(0), A => n13346, ZN => n13344);
   U11795 : OAI22_X1 port map( A1 => n10637, A2 => n261, B1 => n4867, B2 => 
                           n122, ZN => n13346);
   U11796 : AOI22_X1 port map( A1 => n13348, A2 => n4871, B1 => n13349, B2 => 
                           n4873, ZN => n13343);
   U11797 : AOI22_X1 port map( A1 => n13350, A2 => n4875, B1 => n13351, B2 => 
                           n4869, ZN => n13342);
   U11798 : NAND3_X1 port map( A1 => n13352, A2 => n13353, A3 => n13354, ZN => 
                           n11999);
   U11799 : AOI221_X1 port map( B1 => n13345, B2 => n4879, C1 => n171, C2 => 
                           MEM_IN(1), A => n13355, ZN => n13354);
   U11800 : OAI22_X1 port map( A1 => n10636, A2 => n261, B1 => n4881, B2 => 
                           n122, ZN => n13355);
   U11801 : AOI22_X1 port map( A1 => n13348, A2 => n4883, B1 => n13349, B2 => 
                           n4884, ZN => n13353);
   U11802 : AOI22_X1 port map( A1 => n13350, A2 => n4885, B1 => n13351, B2 => 
                           n4882, ZN => n13352);
   U11803 : NAND3_X1 port map( A1 => n13356, A2 => n13357, A3 => n13358, ZN => 
                           n11998);
   U11804 : AOI221_X1 port map( B1 => n13345, B2 => n4889, C1 => n171, C2 => 
                           MEM_IN(2), A => n13359, ZN => n13358);
   U11805 : OAI22_X1 port map( A1 => n10635, A2 => n261, B1 => n4891, B2 => 
                           n122, ZN => n13359);
   U11806 : AOI22_X1 port map( A1 => n13348, A2 => n4893, B1 => n13349, B2 => 
                           n4894, ZN => n13357);
   U11807 : AOI22_X1 port map( A1 => n13350, A2 => n4895, B1 => n13351, B2 => 
                           n4892, ZN => n13356);
   U11808 : NAND3_X1 port map( A1 => n13360, A2 => n13361, A3 => n13362, ZN => 
                           n11997);
   U11809 : AOI221_X1 port map( B1 => n13345, B2 => n4899, C1 => n171, C2 => 
                           MEM_IN(3), A => n13363, ZN => n13362);
   U11810 : OAI22_X1 port map( A1 => n10634, A2 => n261, B1 => n4901, B2 => 
                           n122, ZN => n13363);
   U11811 : AOI22_X1 port map( A1 => n13348, A2 => n4903, B1 => n13349, B2 => 
                           n4904, ZN => n13361);
   U11812 : AOI22_X1 port map( A1 => n13350, A2 => n4905, B1 => n13351, B2 => 
                           n4902, ZN => n13360);
   U11813 : NAND3_X1 port map( A1 => n13364, A2 => n13365, A3 => n13366, ZN => 
                           n11996);
   U11814 : AOI221_X1 port map( B1 => n13345, B2 => n4909, C1 => n171, C2 => 
                           MEM_IN(4), A => n13367, ZN => n13366);
   U11815 : OAI22_X1 port map( A1 => n10633, A2 => n261, B1 => n4911, B2 => 
                           n122, ZN => n13367);
   U11816 : AOI22_X1 port map( A1 => n13348, A2 => n4913, B1 => n13349, B2 => 
                           n4914, ZN => n13365);
   U11817 : AOI22_X1 port map( A1 => n13350, A2 => n4915, B1 => n13351, B2 => 
                           n4912, ZN => n13364);
   U11818 : NAND3_X1 port map( A1 => n13368, A2 => n13369, A3 => n13370, ZN => 
                           n11995);
   U11819 : AOI221_X1 port map( B1 => n13345, B2 => n4919, C1 => n171, C2 => 
                           MEM_IN(5), A => n13371, ZN => n13370);
   U11820 : OAI22_X1 port map( A1 => n10632, A2 => n261, B1 => n4921, B2 => 
                           n122, ZN => n13371);
   U11821 : AOI22_X1 port map( A1 => n13348, A2 => n4923, B1 => n13349, B2 => 
                           n4924, ZN => n13369);
   U11822 : AOI22_X1 port map( A1 => n13350, A2 => n4925, B1 => n13351, B2 => 
                           n4922, ZN => n13368);
   U11823 : NAND3_X1 port map( A1 => n13372, A2 => n13373, A3 => n13374, ZN => 
                           n11994);
   U11824 : AOI221_X1 port map( B1 => n13345, B2 => n4929, C1 => n171, C2 => 
                           MEM_IN(6), A => n13375, ZN => n13374);
   U11825 : OAI22_X1 port map( A1 => n10631, A2 => n261, B1 => n4931, B2 => 
                           n122, ZN => n13375);
   U11826 : AOI22_X1 port map( A1 => n13348, A2 => n4933, B1 => n13349, B2 => 
                           n4934, ZN => n13373);
   U11827 : AOI22_X1 port map( A1 => n13350, A2 => n4935, B1 => n13351, B2 => 
                           n4932, ZN => n13372);
   U11828 : NAND3_X1 port map( A1 => n13376, A2 => n13377, A3 => n13378, ZN => 
                           n11993);
   U11829 : AOI221_X1 port map( B1 => n13345, B2 => n4939, C1 => n171, C2 => 
                           MEM_IN(7), A => n13379, ZN => n13378);
   U11830 : OAI22_X1 port map( A1 => n10630, A2 => n261, B1 => n4941, B2 => 
                           n122, ZN => n13379);
   U11831 : AOI22_X1 port map( A1 => n13348, A2 => n4943, B1 => n13349, B2 => 
                           n4944, ZN => n13377);
   U11832 : AOI22_X1 port map( A1 => n13350, A2 => n4945, B1 => n13351, B2 => 
                           n4942, ZN => n13376);
   U11833 : NAND3_X1 port map( A1 => n13380, A2 => n13381, A3 => n13382, ZN => 
                           n11992);
   U11834 : AOI221_X1 port map( B1 => n13345, B2 => n4949, C1 => n171, C2 => 
                           MEM_IN(8), A => n13383, ZN => n13382);
   U11835 : OAI22_X1 port map( A1 => n10629, A2 => n261, B1 => n4951, B2 => 
                           n122, ZN => n13383);
   U11836 : AOI22_X1 port map( A1 => n13348, A2 => n4953, B1 => n13349, B2 => 
                           n4954, ZN => n13381);
   U11837 : AOI22_X1 port map( A1 => n13350, A2 => n4955, B1 => n13351, B2 => 
                           n4952, ZN => n13380);
   U11838 : NAND3_X1 port map( A1 => n13384, A2 => n13385, A3 => n13386, ZN => 
                           n11991);
   U11839 : AOI221_X1 port map( B1 => n13345, B2 => n4959, C1 => n171, C2 => 
                           MEM_IN(9), A => n13387, ZN => n13386);
   U11840 : OAI22_X1 port map( A1 => n10628, A2 => n261, B1 => n4961, B2 => 
                           n122, ZN => n13387);
   U11841 : AOI22_X1 port map( A1 => n13348, A2 => n4963, B1 => n13349, B2 => 
                           n4964, ZN => n13385);
   U11842 : AOI22_X1 port map( A1 => n13350, A2 => n4965, B1 => n13351, B2 => 
                           n4962, ZN => n13384);
   U11843 : NAND3_X1 port map( A1 => n13388, A2 => n13389, A3 => n13390, ZN => 
                           n11990);
   U11844 : AOI221_X1 port map( B1 => n13345, B2 => n4969, C1 => n171, C2 => 
                           MEM_IN(10), A => n13391, ZN => n13390);
   U11845 : OAI22_X1 port map( A1 => n10627, A2 => n261, B1 => n4971, B2 => 
                           n122, ZN => n13391);
   U11846 : AOI22_X1 port map( A1 => n13348, A2 => n4973, B1 => n13349, B2 => 
                           n4974, ZN => n13389);
   U11847 : AOI22_X1 port map( A1 => n13350, A2 => n4975, B1 => n13351, B2 => 
                           n4972, ZN => n13388);
   U11848 : NAND3_X1 port map( A1 => n13392, A2 => n13393, A3 => n13394, ZN => 
                           n11989);
   U11849 : AOI221_X1 port map( B1 => n13345, B2 => n4979, C1 => n171, C2 => 
                           MEM_IN(11), A => n13395, ZN => n13394);
   U11850 : OAI22_X1 port map( A1 => n10626, A2 => n261, B1 => n4981, B2 => 
                           n122, ZN => n13395);
   U11851 : AOI22_X1 port map( A1 => n13348, A2 => n4983, B1 => n13349, B2 => 
                           n4984, ZN => n13393);
   U11852 : AOI22_X1 port map( A1 => n13350, A2 => n4985, B1 => n13351, B2 => 
                           n4982, ZN => n13392);
   U11853 : NAND3_X1 port map( A1 => n13396, A2 => n13397, A3 => n13398, ZN => 
                           n11988);
   U11854 : AOI221_X1 port map( B1 => n13345, B2 => n4989, C1 => n171, C2 => 
                           MEM_IN(12), A => n13399, ZN => n13398);
   U11855 : OAI22_X1 port map( A1 => n10625, A2 => n261, B1 => n4991, B2 => 
                           n122, ZN => n13399);
   U11856 : AOI22_X1 port map( A1 => n13348, A2 => n4993, B1 => n13349, B2 => 
                           n4994, ZN => n13397);
   U11857 : AOI22_X1 port map( A1 => n13350, A2 => n4995, B1 => n13351, B2 => 
                           n4992, ZN => n13396);
   U11858 : NAND3_X1 port map( A1 => n13400, A2 => n13401, A3 => n13402, ZN => 
                           n11987);
   U11859 : AOI221_X1 port map( B1 => n13345, B2 => n4999, C1 => n171, C2 => 
                           MEM_IN(13), A => n13403, ZN => n13402);
   U11860 : OAI22_X1 port map( A1 => n10624, A2 => n261, B1 => n5001, B2 => 
                           n122, ZN => n13403);
   U11861 : AOI22_X1 port map( A1 => n13348, A2 => n5003, B1 => n13349, B2 => 
                           n5004, ZN => n13401);
   U11862 : AOI22_X1 port map( A1 => n13350, A2 => n5005, B1 => n13351, B2 => 
                           n5002, ZN => n13400);
   U11863 : NAND3_X1 port map( A1 => n13404, A2 => n13405, A3 => n13406, ZN => 
                           n11986);
   U11864 : AOI221_X1 port map( B1 => n13345, B2 => n5009, C1 => n171, C2 => 
                           MEM_IN(14), A => n13407, ZN => n13406);
   U11865 : OAI22_X1 port map( A1 => n10623, A2 => n261, B1 => n5011, B2 => 
                           n122, ZN => n13407);
   U11866 : AOI22_X1 port map( A1 => n13348, A2 => n5013, B1 => n13349, B2 => 
                           n5014, ZN => n13405);
   U11867 : AOI22_X1 port map( A1 => n13350, A2 => n5015, B1 => n13351, B2 => 
                           n5012, ZN => n13404);
   U11868 : NAND3_X1 port map( A1 => n13408, A2 => n13409, A3 => n13410, ZN => 
                           n11985);
   U11869 : AOI221_X1 port map( B1 => n13345, B2 => n5019, C1 => n171, C2 => 
                           MEM_IN(15), A => n13411, ZN => n13410);
   U11870 : OAI22_X1 port map( A1 => n10622, A2 => n261, B1 => n5021, B2 => 
                           n122, ZN => n13411);
   U11871 : AOI22_X1 port map( A1 => n13348, A2 => n5023, B1 => n13349, B2 => 
                           n5024, ZN => n13409);
   U11872 : AOI22_X1 port map( A1 => n13350, A2 => n5025, B1 => n13351, B2 => 
                           n5022, ZN => n13408);
   U11873 : NAND3_X1 port map( A1 => n13412, A2 => n13413, A3 => n13414, ZN => 
                           n11984);
   U11874 : AOI221_X1 port map( B1 => n13345, B2 => n5029, C1 => n171, C2 => 
                           MEM_IN(16), A => n13415, ZN => n13414);
   U11875 : OAI22_X1 port map( A1 => n10621, A2 => n261, B1 => n5031, B2 => 
                           n122, ZN => n13415);
   U11876 : AOI22_X1 port map( A1 => n13348, A2 => n5033, B1 => n13349, B2 => 
                           n5034, ZN => n13413);
   U11877 : AOI22_X1 port map( A1 => n13350, A2 => n5035, B1 => n13351, B2 => 
                           n5032, ZN => n13412);
   U11878 : NAND3_X1 port map( A1 => n13416, A2 => n13417, A3 => n13418, ZN => 
                           n11983);
   U11879 : AOI221_X1 port map( B1 => n13345, B2 => n5039, C1 => n171, C2 => 
                           MEM_IN(17), A => n13419, ZN => n13418);
   U11880 : OAI22_X1 port map( A1 => n10620, A2 => n261, B1 => n5041, B2 => 
                           n122, ZN => n13419);
   U11881 : AOI22_X1 port map( A1 => n13348, A2 => n5043, B1 => n13349, B2 => 
                           n5044, ZN => n13417);
   U11882 : AOI22_X1 port map( A1 => n13350, A2 => n5045, B1 => n13351, B2 => 
                           n5042, ZN => n13416);
   U11883 : NAND3_X1 port map( A1 => n13420, A2 => n13421, A3 => n13422, ZN => 
                           n11982);
   U11884 : AOI221_X1 port map( B1 => n13345, B2 => n5049, C1 => n171, C2 => 
                           MEM_IN(18), A => n13423, ZN => n13422);
   U11885 : OAI22_X1 port map( A1 => n10619, A2 => n261, B1 => n5051, B2 => 
                           n122, ZN => n13423);
   U11886 : AOI22_X1 port map( A1 => n13348, A2 => n5053, B1 => n13349, B2 => 
                           n5054, ZN => n13421);
   U11887 : AOI22_X1 port map( A1 => n13350, A2 => n5055, B1 => n13351, B2 => 
                           n5052, ZN => n13420);
   U11888 : NAND3_X1 port map( A1 => n13424, A2 => n13425, A3 => n13426, ZN => 
                           n11981);
   U11889 : AOI221_X1 port map( B1 => n13345, B2 => n5059, C1 => n171, C2 => 
                           MEM_IN(19), A => n13427, ZN => n13426);
   U11890 : OAI22_X1 port map( A1 => n10618, A2 => n261, B1 => n5061, B2 => 
                           n122, ZN => n13427);
   U11891 : AOI22_X1 port map( A1 => n13348, A2 => n5063, B1 => n13349, B2 => 
                           n5064, ZN => n13425);
   U11892 : AOI22_X1 port map( A1 => n13350, A2 => n5065, B1 => n13351, B2 => 
                           n5062, ZN => n13424);
   U11893 : NAND3_X1 port map( A1 => n13428, A2 => n13429, A3 => n13430, ZN => 
                           n11980);
   U11894 : AOI221_X1 port map( B1 => n13345, B2 => n5069, C1 => n171, C2 => 
                           MEM_IN(20), A => n13431, ZN => n13430);
   U11895 : OAI22_X1 port map( A1 => n10617, A2 => n261, B1 => n5071, B2 => 
                           n122, ZN => n13431);
   U11896 : AOI22_X1 port map( A1 => n13348, A2 => n5073, B1 => n13349, B2 => 
                           n5074, ZN => n13429);
   U11897 : AOI22_X1 port map( A1 => n13350, A2 => n5075, B1 => n13351, B2 => 
                           n5072, ZN => n13428);
   U11898 : NAND3_X1 port map( A1 => n13432, A2 => n13433, A3 => n13434, ZN => 
                           n11979);
   U11899 : AOI221_X1 port map( B1 => n13345, B2 => n5079, C1 => n171, C2 => 
                           MEM_IN(21), A => n13435, ZN => n13434);
   U11900 : OAI22_X1 port map( A1 => n10616, A2 => n261, B1 => n5081, B2 => 
                           n122, ZN => n13435);
   U11901 : AOI22_X1 port map( A1 => n13348, A2 => n5083, B1 => n13349, B2 => 
                           n5084, ZN => n13433);
   U11902 : AOI22_X1 port map( A1 => n13350, A2 => n5085, B1 => n13351, B2 => 
                           n5082, ZN => n13432);
   U11903 : NAND3_X1 port map( A1 => n13436, A2 => n13437, A3 => n13438, ZN => 
                           n11978);
   U11904 : AOI221_X1 port map( B1 => n13345, B2 => n5089, C1 => n171, C2 => 
                           MEM_IN(22), A => n13439, ZN => n13438);
   U11905 : OAI22_X1 port map( A1 => n10615, A2 => n261, B1 => n5091, B2 => 
                           n122, ZN => n13439);
   U11906 : AOI22_X1 port map( A1 => n13348, A2 => n5093, B1 => n13349, B2 => 
                           n5094, ZN => n13437);
   U11907 : AOI22_X1 port map( A1 => n13350, A2 => n5095, B1 => n13351, B2 => 
                           n5092, ZN => n13436);
   U11908 : NAND3_X1 port map( A1 => n13440, A2 => n13441, A3 => n13442, ZN => 
                           n11977);
   U11909 : AOI221_X1 port map( B1 => n13345, B2 => n5099, C1 => n171, C2 => 
                           MEM_IN(23), A => n13443, ZN => n13442);
   U11910 : OAI22_X1 port map( A1 => n10614, A2 => n261, B1 => n5101, B2 => 
                           n122, ZN => n13443);
   U11911 : AOI22_X1 port map( A1 => n13348, A2 => n5103, B1 => n13349, B2 => 
                           n5104, ZN => n13441);
   U11912 : AOI22_X1 port map( A1 => n13350, A2 => n5105, B1 => n13351, B2 => 
                           n5102, ZN => n13440);
   U11913 : NAND3_X1 port map( A1 => n13444, A2 => n13445, A3 => n13446, ZN => 
                           n11976);
   U11914 : AOI221_X1 port map( B1 => n13345, B2 => n5109, C1 => n171, C2 => 
                           MEM_IN(24), A => n13447, ZN => n13446);
   U11915 : OAI22_X1 port map( A1 => n10613, A2 => n261, B1 => n5111, B2 => 
                           n122, ZN => n13447);
   U11916 : AOI22_X1 port map( A1 => n13348, A2 => n5113, B1 => n13349, B2 => 
                           n5114, ZN => n13445);
   U11917 : AOI22_X1 port map( A1 => n13350, A2 => n5115, B1 => n13351, B2 => 
                           n5112, ZN => n13444);
   U11918 : NAND3_X1 port map( A1 => n13448, A2 => n13449, A3 => n13450, ZN => 
                           n11975);
   U11919 : AOI221_X1 port map( B1 => n13345, B2 => n5119, C1 => n171, C2 => 
                           MEM_IN(25), A => n13451, ZN => n13450);
   U11920 : OAI22_X1 port map( A1 => n10612, A2 => n261, B1 => n5121, B2 => 
                           n122, ZN => n13451);
   U11921 : AOI22_X1 port map( A1 => n13348, A2 => n5123, B1 => n13349, B2 => 
                           n5124, ZN => n13449);
   U11922 : AOI22_X1 port map( A1 => n13350, A2 => n5125, B1 => n13351, B2 => 
                           n5122, ZN => n13448);
   U11923 : NAND3_X1 port map( A1 => n13452, A2 => n13453, A3 => n13454, ZN => 
                           n11974);
   U11924 : AOI221_X1 port map( B1 => n13345, B2 => n5129, C1 => n171, C2 => 
                           MEM_IN(26), A => n13455, ZN => n13454);
   U11925 : OAI22_X1 port map( A1 => n10611, A2 => n261, B1 => n5131, B2 => 
                           n122, ZN => n13455);
   U11926 : AOI22_X1 port map( A1 => n13348, A2 => n5133, B1 => n13349, B2 => 
                           n5134, ZN => n13453);
   U11927 : AOI22_X1 port map( A1 => n13350, A2 => n5135, B1 => n13351, B2 => 
                           n5132, ZN => n13452);
   U11928 : NAND3_X1 port map( A1 => n13456, A2 => n13457, A3 => n13458, ZN => 
                           n11973);
   U11929 : AOI221_X1 port map( B1 => n13345, B2 => n5139, C1 => n171, C2 => 
                           MEM_IN(27), A => n13459, ZN => n13458);
   U11930 : OAI22_X1 port map( A1 => n10610, A2 => n261, B1 => n5141, B2 => 
                           n122, ZN => n13459);
   U11931 : AOI22_X1 port map( A1 => n13348, A2 => n5143, B1 => n13349, B2 => 
                           n5144, ZN => n13457);
   U11932 : AOI22_X1 port map( A1 => n13350, A2 => n5145, B1 => n13351, B2 => 
                           n5142, ZN => n13456);
   U11933 : NAND3_X1 port map( A1 => n13460, A2 => n13461, A3 => n13462, ZN => 
                           n11972);
   U11934 : AOI221_X1 port map( B1 => n13345, B2 => n5149, C1 => n171, C2 => 
                           MEM_IN(28), A => n13463, ZN => n13462);
   U11935 : OAI22_X1 port map( A1 => n10609, A2 => n261, B1 => n5151, B2 => 
                           n122, ZN => n13463);
   U11936 : AOI22_X1 port map( A1 => n13348, A2 => n5153, B1 => n13349, B2 => 
                           n5154, ZN => n13461);
   U11937 : AOI22_X1 port map( A1 => n13350, A2 => n5155, B1 => n13351, B2 => 
                           n5152, ZN => n13460);
   U11938 : NAND3_X1 port map( A1 => n13464, A2 => n13465, A3 => n13466, ZN => 
                           n11971);
   U11939 : AOI221_X1 port map( B1 => n13345, B2 => n5159, C1 => n171, C2 => 
                           MEM_IN(29), A => n13467, ZN => n13466);
   U11940 : OAI22_X1 port map( A1 => n10608, A2 => n261, B1 => n5161, B2 => 
                           n122, ZN => n13467);
   U11941 : AOI22_X1 port map( A1 => n13348, A2 => n5163, B1 => n13349, B2 => 
                           n5164, ZN => n13465);
   U11942 : AOI22_X1 port map( A1 => n13350, A2 => n5165, B1 => n13351, B2 => 
                           n5162, ZN => n13464);
   U11943 : NAND3_X1 port map( A1 => n13468, A2 => n13469, A3 => n13470, ZN => 
                           n11970);
   U11944 : AOI221_X1 port map( B1 => n13345, B2 => n5169, C1 => n171, C2 => 
                           MEM_IN(30), A => n13471, ZN => n13470);
   U11945 : OAI22_X1 port map( A1 => n10607, A2 => n261, B1 => n5171, B2 => 
                           n122, ZN => n13471);
   U11946 : AOI22_X1 port map( A1 => n13348, A2 => n5173, B1 => n13349, B2 => 
                           n5174, ZN => n13469);
   U11947 : AOI22_X1 port map( A1 => n13350, A2 => n5175, B1 => n13351, B2 => 
                           n5172, ZN => n13468);
   U11948 : NAND3_X1 port map( A1 => n13472, A2 => n13473, A3 => n13474, ZN => 
                           n11969);
   U11949 : AOI221_X1 port map( B1 => n13345, B2 => n5179, C1 => n171, C2 => 
                           MEM_IN(31), A => n13475, ZN => n13474);
   U11950 : OAI22_X1 port map( A1 => n10606, A2 => n261, B1 => n5181, B2 => 
                           n122, ZN => n13475);
   U11951 : INV_X1 port map( A => n13479, ZN => n13478);
   U11952 : AOI22_X1 port map( A1 => n13348, A2 => n5192, B1 => n13349, B2 => 
                           n5195, ZN => n13473);
   U11953 : NOR2_X1 port map( A1 => n9779, A2 => n4787, ZN => n10220);
   U11954 : AOI22_X1 port map( A1 => n13350, A2 => n5196, B1 => n13351, B2 => 
                           n5191, ZN => n13472);
   U11955 : OAI22_X1 port map( A1 => n13479, A2 => n13477, B1 => n208, B2 => 
                           n260, ZN => n13481);
   U11956 : NAND3_X1 port map( A1 => n208, A2 => n261, A3 => n9630, ZN => 
                           n13477);
   U11957 : INV_X1 port map( A => n13476, ZN => n9630);
   U11958 : OAI22_X1 port map( A1 => n4786, A2 => n13483, B1 => n13484, B2 => 
                           n5204, ZN => n13347);
   U11959 : NOR2_X1 port map( A1 => n13476, A2 => n13479, ZN => n13484);
   U11960 : NAND3_X1 port map( A1 => n10224, A2 => n13485, A3 => n13337, ZN => 
                           n13476);
   U11961 : INV_X1 port map( A => n13486, ZN => n10224);
   U11962 : INV_X1 port map( A => n13487, ZN => n13483);
   U11963 : OAI211_X1 port map( C1 => n13339, C2 => n5923, A => n13480, B => 
                           n5368, ZN => n13487);
   U11964 : AOI21_X1 port map( B1 => n13486, B2 => n5206, A => n13482, ZN => 
                           n13480);
   U11965 : NAND2_X1 port map( A1 => n10072, A2 => n13488, ZN => n13486);
   U11966 : AND2_X1 port map( A1 => n13489, A2 => n9779, ZN => n10072);
   U11967 : NAND2_X1 port map( A1 => n10080, A2 => n5926, ZN => n9779);
   U11968 : NAND3_X1 port map( A1 => n11857, A2 => n10076, A3 => n10225, ZN => 
                           n5923);
   U11969 : NAND3_X1 port map( A1 => n13490, A2 => n11870, A3 => n13491, ZN => 
                           n13479);
   U11970 : NAND3_X1 port map( A1 => n13492, A2 => n13493, A3 => n13494, ZN => 
                           n11968);
   U11971 : AOI221_X1 port map( B1 => n13495, B2 => n4863, C1 => n168, C2 => 
                           MEM_IN(0), A => n13496, ZN => n13494);
   U11972 : OAI22_X1 port map( A1 => n10605, A2 => n245, B1 => n4867, B2 => 
                           n123, ZN => n13496);
   U11973 : AOI22_X1 port map( A1 => n229, A2 => n4873, B1 => n13498, B2 => 
                           n4875, ZN => n13493);
   U11974 : AOI22_X1 port map( A1 => n13499, A2 => n4871, B1 => n13500, B2 => 
                           n4869, ZN => n13492);
   U11975 : NAND3_X1 port map( A1 => n13501, A2 => n13502, A3 => n13503, ZN => 
                           n11967);
   U11976 : AOI221_X1 port map( B1 => n13495, B2 => n4879, C1 => n168, C2 => 
                           MEM_IN(1), A => n13504, ZN => n13503);
   U11977 : OAI22_X1 port map( A1 => n10604, A2 => n245, B1 => n4881, B2 => 
                           n123, ZN => n13504);
   U11978 : AOI22_X1 port map( A1 => n229, A2 => n4884, B1 => n13498, B2 => 
                           n4885, ZN => n13502);
   U11979 : AOI22_X1 port map( A1 => n13499, A2 => n4883, B1 => n13500, B2 => 
                           n4882, ZN => n13501);
   U11980 : NAND3_X1 port map( A1 => n13505, A2 => n13506, A3 => n13507, ZN => 
                           n11966);
   U11981 : AOI221_X1 port map( B1 => n13495, B2 => n4889, C1 => n168, C2 => 
                           MEM_IN(2), A => n13508, ZN => n13507);
   U11982 : OAI22_X1 port map( A1 => n10603, A2 => n245, B1 => n4891, B2 => 
                           n123, ZN => n13508);
   U11983 : AOI22_X1 port map( A1 => n229, A2 => n4894, B1 => n13498, B2 => 
                           n4895, ZN => n13506);
   U11984 : AOI22_X1 port map( A1 => n13499, A2 => n4893, B1 => n13500, B2 => 
                           n4892, ZN => n13505);
   U11985 : NAND3_X1 port map( A1 => n13509, A2 => n13510, A3 => n13511, ZN => 
                           n11965);
   U11986 : AOI221_X1 port map( B1 => n13495, B2 => n4899, C1 => n168, C2 => 
                           MEM_IN(3), A => n13512, ZN => n13511);
   U11987 : OAI22_X1 port map( A1 => n10602, A2 => n245, B1 => n4901, B2 => 
                           n123, ZN => n13512);
   U11988 : AOI22_X1 port map( A1 => n229, A2 => n4904, B1 => n13498, B2 => 
                           n4905, ZN => n13510);
   U11989 : AOI22_X1 port map( A1 => n13499, A2 => n4903, B1 => n13500, B2 => 
                           n4902, ZN => n13509);
   U11990 : NAND3_X1 port map( A1 => n13513, A2 => n13514, A3 => n13515, ZN => 
                           n11964);
   U11991 : AOI221_X1 port map( B1 => n13495, B2 => n4909, C1 => n168, C2 => 
                           MEM_IN(4), A => n13516, ZN => n13515);
   U11992 : OAI22_X1 port map( A1 => n10601, A2 => n245, B1 => n4911, B2 => 
                           n123, ZN => n13516);
   U11993 : AOI22_X1 port map( A1 => n229, A2 => n4914, B1 => n13498, B2 => 
                           n4915, ZN => n13514);
   U11994 : AOI22_X1 port map( A1 => n13499, A2 => n4913, B1 => n13500, B2 => 
                           n4912, ZN => n13513);
   U11995 : NAND3_X1 port map( A1 => n13517, A2 => n13518, A3 => n13519, ZN => 
                           n11963);
   U11996 : AOI221_X1 port map( B1 => n13495, B2 => n4919, C1 => n168, C2 => 
                           MEM_IN(5), A => n13520, ZN => n13519);
   U11997 : OAI22_X1 port map( A1 => n10600, A2 => n245, B1 => n4921, B2 => 
                           n123, ZN => n13520);
   U11998 : AOI22_X1 port map( A1 => n229, A2 => n4924, B1 => n13498, B2 => 
                           n4925, ZN => n13518);
   U11999 : AOI22_X1 port map( A1 => n13499, A2 => n4923, B1 => n13500, B2 => 
                           n4922, ZN => n13517);
   U12000 : NAND3_X1 port map( A1 => n13521, A2 => n13522, A3 => n13523, ZN => 
                           n11962);
   U12001 : AOI221_X1 port map( B1 => n13495, B2 => n4929, C1 => n168, C2 => 
                           MEM_IN(6), A => n13524, ZN => n13523);
   U12002 : OAI22_X1 port map( A1 => n10599, A2 => n245, B1 => n4931, B2 => 
                           n123, ZN => n13524);
   U12003 : AOI22_X1 port map( A1 => n229, A2 => n4934, B1 => n13498, B2 => 
                           n4935, ZN => n13522);
   U12004 : AOI22_X1 port map( A1 => n13499, A2 => n4933, B1 => n13500, B2 => 
                           n4932, ZN => n13521);
   U12005 : NAND3_X1 port map( A1 => n13525, A2 => n13526, A3 => n13527, ZN => 
                           n11961);
   U12006 : AOI221_X1 port map( B1 => n13495, B2 => n4939, C1 => n168, C2 => 
                           MEM_IN(7), A => n13528, ZN => n13527);
   U12007 : OAI22_X1 port map( A1 => n10598, A2 => n245, B1 => n4941, B2 => 
                           n123, ZN => n13528);
   U12008 : AOI22_X1 port map( A1 => n229, A2 => n4944, B1 => n13498, B2 => 
                           n4945, ZN => n13526);
   U12009 : AOI22_X1 port map( A1 => n13499, A2 => n4943, B1 => n13500, B2 => 
                           n4942, ZN => n13525);
   U12010 : NAND3_X1 port map( A1 => n13529, A2 => n13530, A3 => n13531, ZN => 
                           n11960);
   U12011 : AOI221_X1 port map( B1 => n13495, B2 => n4949, C1 => n168, C2 => 
                           MEM_IN(8), A => n13532, ZN => n13531);
   U12012 : OAI22_X1 port map( A1 => n10597, A2 => n245, B1 => n4951, B2 => 
                           n123, ZN => n13532);
   U12013 : AOI22_X1 port map( A1 => n229, A2 => n4954, B1 => n13498, B2 => 
                           n4955, ZN => n13530);
   U12014 : AOI22_X1 port map( A1 => n13499, A2 => n4953, B1 => n13500, B2 => 
                           n4952, ZN => n13529);
   U12015 : NAND3_X1 port map( A1 => n13533, A2 => n13534, A3 => n13535, ZN => 
                           n11959);
   U12016 : AOI221_X1 port map( B1 => n13495, B2 => n4959, C1 => n168, C2 => 
                           MEM_IN(9), A => n13536, ZN => n13535);
   U12017 : OAI22_X1 port map( A1 => n10596, A2 => n245, B1 => n4961, B2 => 
                           n123, ZN => n13536);
   U12018 : AOI22_X1 port map( A1 => n229, A2 => n4964, B1 => n13498, B2 => 
                           n4965, ZN => n13534);
   U12019 : AOI22_X1 port map( A1 => n13499, A2 => n4963, B1 => n13500, B2 => 
                           n4962, ZN => n13533);
   U12020 : NAND3_X1 port map( A1 => n13537, A2 => n13538, A3 => n13539, ZN => 
                           n11958);
   U12021 : AOI221_X1 port map( B1 => n13495, B2 => n4969, C1 => n168, C2 => 
                           MEM_IN(10), A => n13540, ZN => n13539);
   U12022 : OAI22_X1 port map( A1 => n10595, A2 => n245, B1 => n4971, B2 => 
                           n123, ZN => n13540);
   U12023 : AOI22_X1 port map( A1 => n229, A2 => n4974, B1 => n13498, B2 => 
                           n4975, ZN => n13538);
   U12024 : AOI22_X1 port map( A1 => n13499, A2 => n4973, B1 => n13500, B2 => 
                           n4972, ZN => n13537);
   U12025 : NAND3_X1 port map( A1 => n13541, A2 => n13542, A3 => n13543, ZN => 
                           n11957);
   U12026 : AOI221_X1 port map( B1 => n13495, B2 => n4979, C1 => n168, C2 => 
                           MEM_IN(11), A => n13544, ZN => n13543);
   U12027 : OAI22_X1 port map( A1 => n10594, A2 => n245, B1 => n4981, B2 => 
                           n123, ZN => n13544);
   U12028 : AOI22_X1 port map( A1 => n229, A2 => n4984, B1 => n13498, B2 => 
                           n4985, ZN => n13542);
   U12029 : AOI22_X1 port map( A1 => n13499, A2 => n4983, B1 => n13500, B2 => 
                           n4982, ZN => n13541);
   U12030 : NAND3_X1 port map( A1 => n13545, A2 => n13546, A3 => n13547, ZN => 
                           n11956);
   U12031 : AOI221_X1 port map( B1 => n13495, B2 => n4989, C1 => n168, C2 => 
                           MEM_IN(12), A => n13548, ZN => n13547);
   U12032 : OAI22_X1 port map( A1 => n10593, A2 => n245, B1 => n4991, B2 => 
                           n123, ZN => n13548);
   U12033 : AOI22_X1 port map( A1 => n229, A2 => n4994, B1 => n13498, B2 => 
                           n4995, ZN => n13546);
   U12034 : AOI22_X1 port map( A1 => n13499, A2 => n4993, B1 => n13500, B2 => 
                           n4992, ZN => n13545);
   U12035 : NAND3_X1 port map( A1 => n13549, A2 => n13550, A3 => n13551, ZN => 
                           n11955);
   U12036 : AOI221_X1 port map( B1 => n13495, B2 => n4999, C1 => n168, C2 => 
                           MEM_IN(13), A => n13552, ZN => n13551);
   U12037 : OAI22_X1 port map( A1 => n10592, A2 => n245, B1 => n5001, B2 => 
                           n123, ZN => n13552);
   U12038 : AOI22_X1 port map( A1 => n229, A2 => n5004, B1 => n13498, B2 => 
                           n5005, ZN => n13550);
   U12039 : AOI22_X1 port map( A1 => n13499, A2 => n5003, B1 => n13500, B2 => 
                           n5002, ZN => n13549);
   U12040 : NAND3_X1 port map( A1 => n13553, A2 => n13554, A3 => n13555, ZN => 
                           n11954);
   U12041 : AOI221_X1 port map( B1 => n13495, B2 => n5009, C1 => n168, C2 => 
                           MEM_IN(14), A => n13556, ZN => n13555);
   U12042 : OAI22_X1 port map( A1 => n10591, A2 => n245, B1 => n5011, B2 => 
                           n123, ZN => n13556);
   U12043 : AOI22_X1 port map( A1 => n229, A2 => n5014, B1 => n13498, B2 => 
                           n5015, ZN => n13554);
   U12044 : AOI22_X1 port map( A1 => n13499, A2 => n5013, B1 => n13500, B2 => 
                           n5012, ZN => n13553);
   U12045 : NAND3_X1 port map( A1 => n13557, A2 => n13558, A3 => n13559, ZN => 
                           n11953);
   U12046 : AOI221_X1 port map( B1 => n13495, B2 => n5019, C1 => n168, C2 => 
                           MEM_IN(15), A => n13560, ZN => n13559);
   U12047 : OAI22_X1 port map( A1 => n10590, A2 => n245, B1 => n5021, B2 => 
                           n123, ZN => n13560);
   U12048 : AOI22_X1 port map( A1 => n229, A2 => n5024, B1 => n13498, B2 => 
                           n5025, ZN => n13558);
   U12049 : AOI22_X1 port map( A1 => n13499, A2 => n5023, B1 => n13500, B2 => 
                           n5022, ZN => n13557);
   U12050 : NAND3_X1 port map( A1 => n13561, A2 => n13562, A3 => n13563, ZN => 
                           n11952);
   U12051 : AOI221_X1 port map( B1 => n13495, B2 => n5029, C1 => n168, C2 => 
                           MEM_IN(16), A => n13564, ZN => n13563);
   U12052 : OAI22_X1 port map( A1 => n10589, A2 => n245, B1 => n5031, B2 => 
                           n123, ZN => n13564);
   U12053 : AOI22_X1 port map( A1 => n229, A2 => n5034, B1 => n13498, B2 => 
                           n5035, ZN => n13562);
   U12054 : AOI22_X1 port map( A1 => n13499, A2 => n5033, B1 => n13500, B2 => 
                           n5032, ZN => n13561);
   U12055 : NAND3_X1 port map( A1 => n13565, A2 => n13566, A3 => n13567, ZN => 
                           n11951);
   U12056 : AOI221_X1 port map( B1 => n13495, B2 => n5039, C1 => n168, C2 => 
                           MEM_IN(17), A => n13568, ZN => n13567);
   U12057 : OAI22_X1 port map( A1 => n10588, A2 => n245, B1 => n5041, B2 => 
                           n123, ZN => n13568);
   U12058 : AOI22_X1 port map( A1 => n229, A2 => n5044, B1 => n13498, B2 => 
                           n5045, ZN => n13566);
   U12059 : AOI22_X1 port map( A1 => n13499, A2 => n5043, B1 => n13500, B2 => 
                           n5042, ZN => n13565);
   U12060 : NAND3_X1 port map( A1 => n13569, A2 => n13570, A3 => n13571, ZN => 
                           n11950);
   U12061 : AOI221_X1 port map( B1 => n13495, B2 => n5049, C1 => n168, C2 => 
                           MEM_IN(18), A => n13572, ZN => n13571);
   U12062 : OAI22_X1 port map( A1 => n10587, A2 => n245, B1 => n5051, B2 => 
                           n123, ZN => n13572);
   U12063 : AOI22_X1 port map( A1 => n229, A2 => n5054, B1 => n13498, B2 => 
                           n5055, ZN => n13570);
   U12064 : AOI22_X1 port map( A1 => n13499, A2 => n5053, B1 => n13500, B2 => 
                           n5052, ZN => n13569);
   U12065 : NAND3_X1 port map( A1 => n13573, A2 => n13574, A3 => n13575, ZN => 
                           n11949);
   U12066 : AOI221_X1 port map( B1 => n13495, B2 => n5059, C1 => n168, C2 => 
                           MEM_IN(19), A => n13576, ZN => n13575);
   U12067 : OAI22_X1 port map( A1 => n10586, A2 => n245, B1 => n5061, B2 => 
                           n123, ZN => n13576);
   U12068 : AOI22_X1 port map( A1 => n229, A2 => n5064, B1 => n13498, B2 => 
                           n5065, ZN => n13574);
   U12069 : AOI22_X1 port map( A1 => n13499, A2 => n5063, B1 => n13500, B2 => 
                           n5062, ZN => n13573);
   U12070 : NAND3_X1 port map( A1 => n13577, A2 => n13578, A3 => n13579, ZN => 
                           n11948);
   U12071 : AOI221_X1 port map( B1 => n13495, B2 => n5069, C1 => n168, C2 => 
                           MEM_IN(20), A => n13580, ZN => n13579);
   U12072 : OAI22_X1 port map( A1 => n10585, A2 => n245, B1 => n5071, B2 => 
                           n123, ZN => n13580);
   U12073 : AOI22_X1 port map( A1 => n229, A2 => n5074, B1 => n13498, B2 => 
                           n5075, ZN => n13578);
   U12074 : AOI22_X1 port map( A1 => n13499, A2 => n5073, B1 => n13500, B2 => 
                           n5072, ZN => n13577);
   U12075 : NAND3_X1 port map( A1 => n13581, A2 => n13582, A3 => n13583, ZN => 
                           n11947);
   U12076 : AOI221_X1 port map( B1 => n13495, B2 => n5079, C1 => n168, C2 => 
                           MEM_IN(21), A => n13584, ZN => n13583);
   U12077 : OAI22_X1 port map( A1 => n10584, A2 => n245, B1 => n5081, B2 => 
                           n123, ZN => n13584);
   U12078 : AOI22_X1 port map( A1 => n229, A2 => n5084, B1 => n13498, B2 => 
                           n5085, ZN => n13582);
   U12079 : AOI22_X1 port map( A1 => n13499, A2 => n5083, B1 => n13500, B2 => 
                           n5082, ZN => n13581);
   U12080 : NAND3_X1 port map( A1 => n13585, A2 => n13586, A3 => n13587, ZN => 
                           n11946);
   U12081 : AOI221_X1 port map( B1 => n13495, B2 => n5089, C1 => n168, C2 => 
                           MEM_IN(22), A => n13588, ZN => n13587);
   U12082 : OAI22_X1 port map( A1 => n10583, A2 => n245, B1 => n5091, B2 => 
                           n123, ZN => n13588);
   U12083 : AOI22_X1 port map( A1 => n229, A2 => n5094, B1 => n13498, B2 => 
                           n5095, ZN => n13586);
   U12084 : AOI22_X1 port map( A1 => n13499, A2 => n5093, B1 => n13500, B2 => 
                           n5092, ZN => n13585);
   U12085 : NAND3_X1 port map( A1 => n13589, A2 => n13590, A3 => n13591, ZN => 
                           n11945);
   U12086 : AOI221_X1 port map( B1 => n13495, B2 => n5099, C1 => n168, C2 => 
                           MEM_IN(23), A => n13592, ZN => n13591);
   U12087 : OAI22_X1 port map( A1 => n10582, A2 => n245, B1 => n5101, B2 => 
                           n123, ZN => n13592);
   U12088 : AOI22_X1 port map( A1 => n229, A2 => n5104, B1 => n13498, B2 => 
                           n5105, ZN => n13590);
   U12089 : AOI22_X1 port map( A1 => n13499, A2 => n5103, B1 => n13500, B2 => 
                           n5102, ZN => n13589);
   U12090 : NAND3_X1 port map( A1 => n13593, A2 => n13594, A3 => n13595, ZN => 
                           n11944);
   U12091 : AOI221_X1 port map( B1 => n13495, B2 => n5109, C1 => n168, C2 => 
                           MEM_IN(24), A => n13596, ZN => n13595);
   U12092 : OAI22_X1 port map( A1 => n10581, A2 => n245, B1 => n5111, B2 => 
                           n123, ZN => n13596);
   U12093 : AOI22_X1 port map( A1 => n229, A2 => n5114, B1 => n13498, B2 => 
                           n5115, ZN => n13594);
   U12094 : AOI22_X1 port map( A1 => n13499, A2 => n5113, B1 => n13500, B2 => 
                           n5112, ZN => n13593);
   U12095 : NAND3_X1 port map( A1 => n13597, A2 => n13598, A3 => n13599, ZN => 
                           n11943);
   U12096 : AOI221_X1 port map( B1 => n13495, B2 => n5119, C1 => n168, C2 => 
                           MEM_IN(25), A => n13600, ZN => n13599);
   U12097 : OAI22_X1 port map( A1 => n10580, A2 => n245, B1 => n5121, B2 => 
                           n123, ZN => n13600);
   U12098 : AOI22_X1 port map( A1 => n229, A2 => n5124, B1 => n13498, B2 => 
                           n5125, ZN => n13598);
   U12099 : AOI22_X1 port map( A1 => n13499, A2 => n5123, B1 => n13500, B2 => 
                           n5122, ZN => n13597);
   U12100 : NAND3_X1 port map( A1 => n13601, A2 => n13602, A3 => n13603, ZN => 
                           n11942);
   U12101 : AOI221_X1 port map( B1 => n13495, B2 => n5129, C1 => n168, C2 => 
                           MEM_IN(26), A => n13604, ZN => n13603);
   U12102 : OAI22_X1 port map( A1 => n10579, A2 => n245, B1 => n5131, B2 => 
                           n123, ZN => n13604);
   U12103 : AOI22_X1 port map( A1 => n229, A2 => n5134, B1 => n13498, B2 => 
                           n5135, ZN => n13602);
   U12104 : AOI22_X1 port map( A1 => n13499, A2 => n5133, B1 => n13500, B2 => 
                           n5132, ZN => n13601);
   U12105 : NAND3_X1 port map( A1 => n13605, A2 => n13606, A3 => n13607, ZN => 
                           n11941);
   U12106 : AOI221_X1 port map( B1 => n13495, B2 => n5139, C1 => n168, C2 => 
                           MEM_IN(27), A => n13608, ZN => n13607);
   U12107 : OAI22_X1 port map( A1 => n10578, A2 => n245, B1 => n5141, B2 => 
                           n123, ZN => n13608);
   U12108 : AOI22_X1 port map( A1 => n229, A2 => n5144, B1 => n13498, B2 => 
                           n5145, ZN => n13606);
   U12109 : AOI22_X1 port map( A1 => n13499, A2 => n5143, B1 => n13500, B2 => 
                           n5142, ZN => n13605);
   U12110 : NAND3_X1 port map( A1 => n13609, A2 => n13610, A3 => n13611, ZN => 
                           n11940);
   U12111 : AOI221_X1 port map( B1 => n13495, B2 => n5149, C1 => n168, C2 => 
                           MEM_IN(28), A => n13612, ZN => n13611);
   U12112 : OAI22_X1 port map( A1 => n10577, A2 => n245, B1 => n5151, B2 => 
                           n123, ZN => n13612);
   U12113 : AOI22_X1 port map( A1 => n229, A2 => n5154, B1 => n13498, B2 => 
                           n5155, ZN => n13610);
   U12114 : AOI22_X1 port map( A1 => n13499, A2 => n5153, B1 => n13500, B2 => 
                           n5152, ZN => n13609);
   U12115 : NAND3_X1 port map( A1 => n13613, A2 => n13614, A3 => n13615, ZN => 
                           n11939);
   U12116 : AOI221_X1 port map( B1 => n13495, B2 => n5159, C1 => n168, C2 => 
                           MEM_IN(29), A => n13616, ZN => n13615);
   U12117 : OAI22_X1 port map( A1 => n10576, A2 => n245, B1 => n5161, B2 => 
                           n123, ZN => n13616);
   U12118 : AOI22_X1 port map( A1 => n229, A2 => n5164, B1 => n13498, B2 => 
                           n5165, ZN => n13614);
   U12119 : AOI22_X1 port map( A1 => n13499, A2 => n5163, B1 => n13500, B2 => 
                           n5162, ZN => n13613);
   U12120 : NAND3_X1 port map( A1 => n13617, A2 => n13618, A3 => n13619, ZN => 
                           n11938);
   U12121 : AOI221_X1 port map( B1 => n13495, B2 => n5169, C1 => n168, C2 => 
                           MEM_IN(30), A => n13620, ZN => n13619);
   U12122 : OAI22_X1 port map( A1 => n10575, A2 => n245, B1 => n5171, B2 => 
                           n123, ZN => n13620);
   U12123 : AOI22_X1 port map( A1 => n229, A2 => n5174, B1 => n13498, B2 => 
                           n5175, ZN => n13618);
   U12124 : AOI22_X1 port map( A1 => n13499, A2 => n5173, B1 => n13500, B2 => 
                           n5172, ZN => n13617);
   U12125 : NAND3_X1 port map( A1 => n13621, A2 => n13622, A3 => n13623, ZN => 
                           n11937);
   U12126 : AOI221_X1 port map( B1 => n13495, B2 => n5179, C1 => n168, C2 => 
                           MEM_IN(31), A => n13624, ZN => n13623);
   U12127 : OAI22_X1 port map( A1 => n10574, A2 => n245, B1 => n5181, B2 => 
                           n123, ZN => n13624);
   U12128 : INV_X1 port map( A => n13333, ZN => n11849);
   U12129 : AOI22_X1 port map( A1 => n229, A2 => n5195, B1 => n13498, B2 => 
                           n5196, ZN => n13622);
   U12130 : AOI22_X1 port map( A1 => n13499, A2 => n5192, B1 => n13500, B2 => 
                           n5191, ZN => n13621);
   U12131 : INV_X1 port map( A => n13631, ZN => n13629);
   U12132 : AOI22_X1 port map( A1 => n13627, A2 => n13634, B1 => n4841, B2 => 
                           n245, ZN => n13631);
   U12133 : INV_X1 port map( A => n13626, ZN => n13634);
   U12134 : NAND3_X1 port map( A1 => n208, A2 => n245, A3 => n9778, ZN => 
                           n13626);
   U12135 : OAI22_X1 port map( A1 => n4786, A2 => n13635, B1 => n13636, B2 => 
                           n5204, ZN => n13497);
   U12136 : NOR2_X1 port map( A1 => n13625, A2 => n13637, ZN => n13636);
   U12137 : INV_X1 port map( A => n9778, ZN => n13625);
   U12138 : NOR3_X1 port map( A1 => n10079, A2 => n9928, A3 => n13638, ZN => 
                           n9778);
   U12139 : INV_X1 port map( A => n13489, ZN => n9928);
   U12140 : AOI211_X1 port map( C1 => n10073, C2 => n8448, A => n13639, B => 
                           n13333, ZN => n13635);
   U12141 : NOR2_X1 port map( A1 => n13489, A2 => n4787, ZN => n13333);
   U12142 : NAND2_X1 port map( A1 => n10080, A2 => n6079, ZN => n13489);
   U12143 : INV_X1 port map( A => n6076, ZN => n8448);
   U12144 : NAND3_X1 port map( A1 => n10076, A2 => n10077, A3 => n11857, ZN => 
                           n6076);
   U12145 : INV_X1 port map( A => n13637, ZN => n13627);
   U12146 : NAND2_X1 port map( A1 => n13640, A2 => n11870, ZN => n13637);
   U12147 : OAI21_X1 port map( B1 => n13641, B2 => n13642, A => n10226, ZN => 
                           n11870);
   U12148 : INV_X1 port map( A => n13643, ZN => n13641);
   U12149 : NAND3_X1 port map( A1 => n13644, A2 => n13645, A3 => n13646, ZN => 
                           n11936);
   U12150 : AOI221_X1 port map( B1 => n13647, B2 => n4863, C1 => n13648, C2 => 
                           MEM_IN(0), A => n13649, ZN => n13646);
   U12151 : OAI22_X1 port map( A1 => n10573, A2 => n249, B1 => n4867, B2 => 
                           n120, ZN => n13649);
   U12152 : AOI22_X1 port map( A1 => n13651, A2 => n4873, B1 => n153, B2 => 
                           n4869, ZN => n13645);
   U12153 : AOI22_X1 port map( A1 => n13652, A2 => n4875, B1 => n13653, B2 => 
                           n4871, ZN => n13644);
   U12154 : NAND3_X1 port map( A1 => n13654, A2 => n13655, A3 => n13656, ZN => 
                           n11935);
   U12155 : AOI221_X1 port map( B1 => n13647, B2 => n4879, C1 => n13648, C2 => 
                           MEM_IN(1), A => n13657, ZN => n13656);
   U12156 : OAI22_X1 port map( A1 => n10572, A2 => n249, B1 => n4881, B2 => 
                           n120, ZN => n13657);
   U12157 : AOI22_X1 port map( A1 => n13651, A2 => n4884, B1 => n153, B2 => 
                           n4882, ZN => n13655);
   U12158 : AOI22_X1 port map( A1 => n13652, A2 => n4885, B1 => n13653, B2 => 
                           n4883, ZN => n13654);
   U12159 : NAND3_X1 port map( A1 => n13658, A2 => n13659, A3 => n13660, ZN => 
                           n11934);
   U12160 : AOI221_X1 port map( B1 => n13647, B2 => n4889, C1 => n13648, C2 => 
                           MEM_IN(2), A => n13661, ZN => n13660);
   U12161 : OAI22_X1 port map( A1 => n10571, A2 => n249, B1 => n4891, B2 => 
                           n120, ZN => n13661);
   U12162 : AOI22_X1 port map( A1 => n13651, A2 => n4894, B1 => n153, B2 => 
                           n4892, ZN => n13659);
   U12163 : AOI22_X1 port map( A1 => n13652, A2 => n4895, B1 => n13653, B2 => 
                           n4893, ZN => n13658);
   U12164 : NAND3_X1 port map( A1 => n13662, A2 => n13663, A3 => n13664, ZN => 
                           n11933);
   U12165 : AOI221_X1 port map( B1 => n13647, B2 => n4899, C1 => n13648, C2 => 
                           MEM_IN(3), A => n13665, ZN => n13664);
   U12166 : OAI22_X1 port map( A1 => n10570, A2 => n249, B1 => n4901, B2 => 
                           n120, ZN => n13665);
   U12167 : AOI22_X1 port map( A1 => n13651, A2 => n4904, B1 => n153, B2 => 
                           n4902, ZN => n13663);
   U12168 : AOI22_X1 port map( A1 => n13652, A2 => n4905, B1 => n13653, B2 => 
                           n4903, ZN => n13662);
   U12169 : NAND3_X1 port map( A1 => n13666, A2 => n13667, A3 => n13668, ZN => 
                           n11932);
   U12170 : AOI221_X1 port map( B1 => n13647, B2 => n4909, C1 => n13648, C2 => 
                           MEM_IN(4), A => n13669, ZN => n13668);
   U12171 : OAI22_X1 port map( A1 => n10569, A2 => n249, B1 => n4911, B2 => 
                           n120, ZN => n13669);
   U12172 : AOI22_X1 port map( A1 => n13651, A2 => n4914, B1 => n153, B2 => 
                           n4912, ZN => n13667);
   U12173 : AOI22_X1 port map( A1 => n13652, A2 => n4915, B1 => n13653, B2 => 
                           n4913, ZN => n13666);
   U12174 : NAND3_X1 port map( A1 => n13670, A2 => n13671, A3 => n13672, ZN => 
                           n11931);
   U12175 : AOI221_X1 port map( B1 => n13647, B2 => n4919, C1 => n13648, C2 => 
                           MEM_IN(5), A => n13673, ZN => n13672);
   U12176 : OAI22_X1 port map( A1 => n10568, A2 => n249, B1 => n4921, B2 => 
                           n120, ZN => n13673);
   U12177 : AOI22_X1 port map( A1 => n13651, A2 => n4924, B1 => n153, B2 => 
                           n4922, ZN => n13671);
   U12178 : AOI22_X1 port map( A1 => n13652, A2 => n4925, B1 => n13653, B2 => 
                           n4923, ZN => n13670);
   U12179 : NAND3_X1 port map( A1 => n13674, A2 => n13675, A3 => n13676, ZN => 
                           n11930);
   U12180 : AOI221_X1 port map( B1 => n13647, B2 => n4929, C1 => n13648, C2 => 
                           MEM_IN(6), A => n13677, ZN => n13676);
   U12181 : OAI22_X1 port map( A1 => n10567, A2 => n249, B1 => n4931, B2 => 
                           n120, ZN => n13677);
   U12182 : AOI22_X1 port map( A1 => n13651, A2 => n4934, B1 => n153, B2 => 
                           n4932, ZN => n13675);
   U12183 : AOI22_X1 port map( A1 => n13652, A2 => n4935, B1 => n13653, B2 => 
                           n4933, ZN => n13674);
   U12184 : NAND3_X1 port map( A1 => n13678, A2 => n13679, A3 => n13680, ZN => 
                           n11929);
   U12185 : AOI221_X1 port map( B1 => n13647, B2 => n4939, C1 => n13648, C2 => 
                           MEM_IN(7), A => n13681, ZN => n13680);
   U12186 : OAI22_X1 port map( A1 => n10566, A2 => n249, B1 => n4941, B2 => 
                           n120, ZN => n13681);
   U12187 : AOI22_X1 port map( A1 => n13651, A2 => n4944, B1 => n153, B2 => 
                           n4942, ZN => n13679);
   U12188 : AOI22_X1 port map( A1 => n13652, A2 => n4945, B1 => n13653, B2 => 
                           n4943, ZN => n13678);
   U12189 : NAND3_X1 port map( A1 => n13682, A2 => n13683, A3 => n13684, ZN => 
                           n11928);
   U12190 : AOI221_X1 port map( B1 => n13647, B2 => n4949, C1 => n13648, C2 => 
                           MEM_IN(8), A => n13685, ZN => n13684);
   U12191 : OAI22_X1 port map( A1 => n10565, A2 => n249, B1 => n4951, B2 => 
                           n120, ZN => n13685);
   U12192 : AOI22_X1 port map( A1 => n13651, A2 => n4954, B1 => n153, B2 => 
                           n4952, ZN => n13683);
   U12193 : AOI22_X1 port map( A1 => n13652, A2 => n4955, B1 => n13653, B2 => 
                           n4953, ZN => n13682);
   U12194 : NAND3_X1 port map( A1 => n13686, A2 => n13687, A3 => n13688, ZN => 
                           n11927);
   U12195 : AOI221_X1 port map( B1 => n13647, B2 => n4959, C1 => n13648, C2 => 
                           MEM_IN(9), A => n13689, ZN => n13688);
   U12196 : OAI22_X1 port map( A1 => n10564, A2 => n249, B1 => n4961, B2 => 
                           n120, ZN => n13689);
   U12197 : AOI22_X1 port map( A1 => n13651, A2 => n4964, B1 => n153, B2 => 
                           n4962, ZN => n13687);
   U12198 : AOI22_X1 port map( A1 => n13652, A2 => n4965, B1 => n13653, B2 => 
                           n4963, ZN => n13686);
   U12199 : NAND3_X1 port map( A1 => n13690, A2 => n13691, A3 => n13692, ZN => 
                           n11926);
   U12200 : AOI221_X1 port map( B1 => n13647, B2 => n4969, C1 => n13648, C2 => 
                           MEM_IN(10), A => n13693, ZN => n13692);
   U12201 : OAI22_X1 port map( A1 => n10563, A2 => n249, B1 => n4971, B2 => 
                           n120, ZN => n13693);
   U12202 : AOI22_X1 port map( A1 => n13651, A2 => n4974, B1 => n153, B2 => 
                           n4972, ZN => n13691);
   U12203 : AOI22_X1 port map( A1 => n13652, A2 => n4975, B1 => n13653, B2 => 
                           n4973, ZN => n13690);
   U12204 : NAND3_X1 port map( A1 => n13694, A2 => n13695, A3 => n13696, ZN => 
                           n11925);
   U12205 : AOI221_X1 port map( B1 => n13647, B2 => n4979, C1 => n13648, C2 => 
                           MEM_IN(11), A => n13697, ZN => n13696);
   U12206 : OAI22_X1 port map( A1 => n10562, A2 => n249, B1 => n4981, B2 => 
                           n120, ZN => n13697);
   U12207 : AOI22_X1 port map( A1 => n13651, A2 => n4984, B1 => n153, B2 => 
                           n4982, ZN => n13695);
   U12208 : AOI22_X1 port map( A1 => n13652, A2 => n4985, B1 => n13653, B2 => 
                           n4983, ZN => n13694);
   U12209 : NAND3_X1 port map( A1 => n13698, A2 => n13699, A3 => n13700, ZN => 
                           n11924);
   U12210 : AOI221_X1 port map( B1 => n13647, B2 => n4989, C1 => n13648, C2 => 
                           MEM_IN(12), A => n13701, ZN => n13700);
   U12211 : OAI22_X1 port map( A1 => n10561, A2 => n249, B1 => n4991, B2 => 
                           n120, ZN => n13701);
   U12212 : AOI22_X1 port map( A1 => n13651, A2 => n4994, B1 => n153, B2 => 
                           n4992, ZN => n13699);
   U12213 : AOI22_X1 port map( A1 => n13652, A2 => n4995, B1 => n13653, B2 => 
                           n4993, ZN => n13698);
   U12214 : NAND3_X1 port map( A1 => n13702, A2 => n13703, A3 => n13704, ZN => 
                           n11923);
   U12215 : AOI221_X1 port map( B1 => n13647, B2 => n4999, C1 => n13648, C2 => 
                           MEM_IN(13), A => n13705, ZN => n13704);
   U12216 : OAI22_X1 port map( A1 => n10560, A2 => n249, B1 => n5001, B2 => 
                           n120, ZN => n13705);
   U12217 : AOI22_X1 port map( A1 => n13651, A2 => n5004, B1 => n153, B2 => 
                           n5002, ZN => n13703);
   U12218 : AOI22_X1 port map( A1 => n13652, A2 => n5005, B1 => n13653, B2 => 
                           n5003, ZN => n13702);
   U12219 : NAND3_X1 port map( A1 => n13706, A2 => n13707, A3 => n13708, ZN => 
                           n11922);
   U12220 : AOI221_X1 port map( B1 => n13647, B2 => n5009, C1 => n13648, C2 => 
                           MEM_IN(14), A => n13709, ZN => n13708);
   U12221 : OAI22_X1 port map( A1 => n10559, A2 => n249, B1 => n5011, B2 => 
                           n120, ZN => n13709);
   U12222 : AOI22_X1 port map( A1 => n13651, A2 => n5014, B1 => n153, B2 => 
                           n5012, ZN => n13707);
   U12223 : AOI22_X1 port map( A1 => n13652, A2 => n5015, B1 => n13653, B2 => 
                           n5013, ZN => n13706);
   U12224 : NAND3_X1 port map( A1 => n13710, A2 => n13711, A3 => n13712, ZN => 
                           n11921);
   U12225 : AOI221_X1 port map( B1 => n13647, B2 => n5019, C1 => n13648, C2 => 
                           MEM_IN(15), A => n13713, ZN => n13712);
   U12226 : OAI22_X1 port map( A1 => n10558, A2 => n249, B1 => n5021, B2 => 
                           n120, ZN => n13713);
   U12227 : AOI22_X1 port map( A1 => n13651, A2 => n5024, B1 => n153, B2 => 
                           n5022, ZN => n13711);
   U12228 : AOI22_X1 port map( A1 => n13652, A2 => n5025, B1 => n13653, B2 => 
                           n5023, ZN => n13710);
   U12229 : NAND3_X1 port map( A1 => n13714, A2 => n13715, A3 => n13716, ZN => 
                           n11920);
   U12230 : AOI221_X1 port map( B1 => n13647, B2 => n5029, C1 => n13648, C2 => 
                           MEM_IN(16), A => n13717, ZN => n13716);
   U12231 : OAI22_X1 port map( A1 => n10557, A2 => n249, B1 => n5031, B2 => 
                           n120, ZN => n13717);
   U12232 : AOI22_X1 port map( A1 => n13651, A2 => n5034, B1 => n153, B2 => 
                           n5032, ZN => n13715);
   U12233 : AOI22_X1 port map( A1 => n13652, A2 => n5035, B1 => n13653, B2 => 
                           n5033, ZN => n13714);
   U12234 : NAND3_X1 port map( A1 => n13718, A2 => n13719, A3 => n13720, ZN => 
                           n11919);
   U12235 : AOI221_X1 port map( B1 => n13647, B2 => n5039, C1 => n13648, C2 => 
                           MEM_IN(17), A => n13721, ZN => n13720);
   U12236 : OAI22_X1 port map( A1 => n10556, A2 => n249, B1 => n5041, B2 => 
                           n120, ZN => n13721);
   U12237 : AOI22_X1 port map( A1 => n13651, A2 => n5044, B1 => n153, B2 => 
                           n5042, ZN => n13719);
   U12238 : AOI22_X1 port map( A1 => n13652, A2 => n5045, B1 => n13653, B2 => 
                           n5043, ZN => n13718);
   U12239 : NAND3_X1 port map( A1 => n13722, A2 => n13723, A3 => n13724, ZN => 
                           n11918);
   U12240 : AOI221_X1 port map( B1 => n13647, B2 => n5049, C1 => n13648, C2 => 
                           MEM_IN(18), A => n13725, ZN => n13724);
   U12241 : OAI22_X1 port map( A1 => n10555, A2 => n249, B1 => n5051, B2 => 
                           n120, ZN => n13725);
   U12242 : AOI22_X1 port map( A1 => n13651, A2 => n5054, B1 => n153, B2 => 
                           n5052, ZN => n13723);
   U12243 : AOI22_X1 port map( A1 => n13652, A2 => n5055, B1 => n13653, B2 => 
                           n5053, ZN => n13722);
   U12244 : NAND3_X1 port map( A1 => n13726, A2 => n13727, A3 => n13728, ZN => 
                           n11917);
   U12245 : AOI221_X1 port map( B1 => n13647, B2 => n5059, C1 => n13648, C2 => 
                           MEM_IN(19), A => n13729, ZN => n13728);
   U12246 : OAI22_X1 port map( A1 => n10554, A2 => n249, B1 => n5061, B2 => 
                           n120, ZN => n13729);
   U12247 : AOI22_X1 port map( A1 => n13651, A2 => n5064, B1 => n153, B2 => 
                           n5062, ZN => n13727);
   U12248 : AOI22_X1 port map( A1 => n13652, A2 => n5065, B1 => n13653, B2 => 
                           n5063, ZN => n13726);
   U12249 : NAND3_X1 port map( A1 => n13730, A2 => n13731, A3 => n13732, ZN => 
                           n11916);
   U12250 : AOI221_X1 port map( B1 => n13647, B2 => n5069, C1 => n13648, C2 => 
                           MEM_IN(20), A => n13733, ZN => n13732);
   U12251 : OAI22_X1 port map( A1 => n10553, A2 => n249, B1 => n5071, B2 => 
                           n120, ZN => n13733);
   U12252 : AOI22_X1 port map( A1 => n13651, A2 => n5074, B1 => n153, B2 => 
                           n5072, ZN => n13731);
   U12253 : AOI22_X1 port map( A1 => n13652, A2 => n5075, B1 => n13653, B2 => 
                           n5073, ZN => n13730);
   U12254 : NAND3_X1 port map( A1 => n13734, A2 => n13735, A3 => n13736, ZN => 
                           n11915);
   U12255 : AOI221_X1 port map( B1 => n13647, B2 => n5079, C1 => n13648, C2 => 
                           MEM_IN(21), A => n13737, ZN => n13736);
   U12256 : OAI22_X1 port map( A1 => n10552, A2 => n249, B1 => n5081, B2 => 
                           n120, ZN => n13737);
   U12257 : AOI22_X1 port map( A1 => n13651, A2 => n5084, B1 => n153, B2 => 
                           n5082, ZN => n13735);
   U12258 : AOI22_X1 port map( A1 => n13652, A2 => n5085, B1 => n13653, B2 => 
                           n5083, ZN => n13734);
   U12259 : NAND3_X1 port map( A1 => n13738, A2 => n13739, A3 => n13740, ZN => 
                           n11914);
   U12260 : AOI221_X1 port map( B1 => n13647, B2 => n5089, C1 => n13648, C2 => 
                           MEM_IN(22), A => n13741, ZN => n13740);
   U12261 : OAI22_X1 port map( A1 => n10551, A2 => n249, B1 => n5091, B2 => 
                           n120, ZN => n13741);
   U12262 : AOI22_X1 port map( A1 => n13651, A2 => n5094, B1 => n153, B2 => 
                           n5092, ZN => n13739);
   U12263 : AOI22_X1 port map( A1 => n13652, A2 => n5095, B1 => n13653, B2 => 
                           n5093, ZN => n13738);
   U12264 : NAND3_X1 port map( A1 => n13742, A2 => n13743, A3 => n13744, ZN => 
                           n11913);
   U12265 : AOI221_X1 port map( B1 => n13647, B2 => n5099, C1 => n13648, C2 => 
                           MEM_IN(23), A => n13745, ZN => n13744);
   U12266 : OAI22_X1 port map( A1 => n10550, A2 => n249, B1 => n5101, B2 => 
                           n120, ZN => n13745);
   U12267 : AOI22_X1 port map( A1 => n13651, A2 => n5104, B1 => n153, B2 => 
                           n5102, ZN => n13743);
   U12268 : AOI22_X1 port map( A1 => n13652, A2 => n5105, B1 => n13653, B2 => 
                           n5103, ZN => n13742);
   U12269 : NAND3_X1 port map( A1 => n13746, A2 => n13747, A3 => n13748, ZN => 
                           n11912);
   U12270 : AOI221_X1 port map( B1 => n13647, B2 => n5109, C1 => n13648, C2 => 
                           MEM_IN(24), A => n13749, ZN => n13748);
   U12271 : OAI22_X1 port map( A1 => n10549, A2 => n249, B1 => n5111, B2 => 
                           n120, ZN => n13749);
   U12272 : AOI22_X1 port map( A1 => n13651, A2 => n5114, B1 => n153, B2 => 
                           n5112, ZN => n13747);
   U12273 : AOI22_X1 port map( A1 => n13652, A2 => n5115, B1 => n13653, B2 => 
                           n5113, ZN => n13746);
   U12274 : NAND3_X1 port map( A1 => n13750, A2 => n13751, A3 => n13752, ZN => 
                           n11911);
   U12275 : AOI221_X1 port map( B1 => n13647, B2 => n5119, C1 => n13648, C2 => 
                           MEM_IN(25), A => n13753, ZN => n13752);
   U12276 : OAI22_X1 port map( A1 => n10548, A2 => n249, B1 => n5121, B2 => 
                           n120, ZN => n13753);
   U12277 : AOI22_X1 port map( A1 => n13651, A2 => n5124, B1 => n153, B2 => 
                           n5122, ZN => n13751);
   U12278 : AOI22_X1 port map( A1 => n13652, A2 => n5125, B1 => n13653, B2 => 
                           n5123, ZN => n13750);
   U12279 : NAND3_X1 port map( A1 => n13754, A2 => n13755, A3 => n13756, ZN => 
                           n11910);
   U12280 : AOI221_X1 port map( B1 => n13647, B2 => n5129, C1 => n13648, C2 => 
                           MEM_IN(26), A => n13757, ZN => n13756);
   U12281 : OAI22_X1 port map( A1 => n10547, A2 => n249, B1 => n5131, B2 => 
                           n120, ZN => n13757);
   U12282 : AOI22_X1 port map( A1 => n13651, A2 => n5134, B1 => n153, B2 => 
                           n5132, ZN => n13755);
   U12283 : AOI22_X1 port map( A1 => n13652, A2 => n5135, B1 => n13653, B2 => 
                           n5133, ZN => n13754);
   U12284 : NAND3_X1 port map( A1 => n13758, A2 => n13759, A3 => n13760, ZN => 
                           n11909);
   U12285 : AOI221_X1 port map( B1 => n13647, B2 => n5139, C1 => n13648, C2 => 
                           MEM_IN(27), A => n13761, ZN => n13760);
   U12286 : OAI22_X1 port map( A1 => n10546, A2 => n249, B1 => n5141, B2 => 
                           n120, ZN => n13761);
   U12287 : AOI22_X1 port map( A1 => n13651, A2 => n5144, B1 => n153, B2 => 
                           n5142, ZN => n13759);
   U12288 : AOI22_X1 port map( A1 => n13652, A2 => n5145, B1 => n13653, B2 => 
                           n5143, ZN => n13758);
   U12289 : NAND3_X1 port map( A1 => n13762, A2 => n13763, A3 => n13764, ZN => 
                           n11908);
   U12290 : AOI221_X1 port map( B1 => n13647, B2 => n5149, C1 => n13648, C2 => 
                           MEM_IN(28), A => n13765, ZN => n13764);
   U12291 : OAI22_X1 port map( A1 => n10545, A2 => n249, B1 => n5151, B2 => 
                           n120, ZN => n13765);
   U12292 : AOI22_X1 port map( A1 => n13651, A2 => n5154, B1 => n153, B2 => 
                           n5152, ZN => n13763);
   U12293 : AOI22_X1 port map( A1 => n13652, A2 => n5155, B1 => n13653, B2 => 
                           n5153, ZN => n13762);
   U12294 : NAND3_X1 port map( A1 => n13766, A2 => n13767, A3 => n13768, ZN => 
                           n11907);
   U12295 : AOI221_X1 port map( B1 => n13647, B2 => n5159, C1 => n13648, C2 => 
                           MEM_IN(29), A => n13769, ZN => n13768);
   U12296 : OAI22_X1 port map( A1 => n10544, A2 => n249, B1 => n5161, B2 => 
                           n120, ZN => n13769);
   U12297 : AOI22_X1 port map( A1 => n13651, A2 => n5164, B1 => n153, B2 => 
                           n5162, ZN => n13767);
   U12298 : AOI22_X1 port map( A1 => n13652, A2 => n5165, B1 => n13653, B2 => 
                           n5163, ZN => n13766);
   U12299 : NAND3_X1 port map( A1 => n13770, A2 => n13771, A3 => n13772, ZN => 
                           n11906);
   U12300 : AOI221_X1 port map( B1 => n13647, B2 => n5169, C1 => n13648, C2 => 
                           MEM_IN(30), A => n13773, ZN => n13772);
   U12301 : OAI22_X1 port map( A1 => n10543, A2 => n249, B1 => n5171, B2 => 
                           n120, ZN => n13773);
   U12302 : AOI22_X1 port map( A1 => n13651, A2 => n5174, B1 => n153, B2 => 
                           n5172, ZN => n13771);
   U12303 : AOI22_X1 port map( A1 => n13652, A2 => n5175, B1 => n13653, B2 => 
                           n5173, ZN => n13770);
   U12304 : NAND3_X1 port map( A1 => n13774, A2 => n13775, A3 => n13776, ZN => 
                           n11905);
   U12305 : AOI221_X1 port map( B1 => n13647, B2 => n5179, C1 => n13648, C2 => 
                           MEM_IN(31), A => n13777, ZN => n13776);
   U12306 : OAI22_X1 port map( A1 => n10542, A2 => n249, B1 => n5181, B2 => 
                           n120, ZN => n13777);
   U12307 : AOI22_X1 port map( A1 => n13651, A2 => n5195, B1 => n153, B2 => 
                           n5191, ZN => n13775);
   U12308 : NOR2_X1 port map( A1 => n13632, A2 => n13488, ZN => n13630);
   U12309 : AOI22_X1 port map( A1 => n13652, A2 => n5196, B1 => n13653, B2 => 
                           n5192, ZN => n13774);
   U12310 : INV_X1 port map( A => n13782, ZN => n13780);
   U12311 : AOI22_X1 port map( A1 => n13783, A2 => n13778, B1 => n4841, B2 => 
                           n249, ZN => n13782);
   U12312 : AND3_X1 port map( A1 => n208, A2 => n249, A3 => n13784, ZN => 
                           n13778);
   U12313 : OAI22_X1 port map( A1 => n4786, A2 => n13785, B1 => n13786, B2 => 
                           n5204, ZN => n13650);
   U12314 : NOR2_X1 port map( A1 => n9927, A2 => n13779, ZN => n13786);
   U12315 : INV_X1 port map( A => n13783, ZN => n13779);
   U12316 : INV_X1 port map( A => n13784, ZN => n9927);
   U12317 : AOI211_X1 port map( C1 => n5775, C2 => n10226, A => n10079, B => 
                           n13638, ZN => n13784);
   U12318 : INV_X1 port map( A => n13488, ZN => n10079);
   U12319 : AOI211_X1 port map( C1 => n10073, C2 => n6223, A => n13639, B => 
                           n13787, ZN => n13785);
   U12320 : OAI211_X1 port map( C1 => n13337, C2 => n4787, A => n13331, B => 
                           n5368, ZN => n13639);
   U12321 : INV_X1 port map( A => n13334, ZN => n13331);
   U12322 : NOR2_X1 port map( A1 => n13488, A2 => n4787, ZN => n13334);
   U12323 : NAND2_X1 port map( A1 => n10080, A2 => n6228, ZN => n13488);
   U12324 : INV_X1 port map( A => n8594, ZN => n6223);
   U12325 : NAND3_X1 port map( A1 => n10075, A2 => n10076, A3 => n10225, ZN => 
                           n8594);
   U12326 : AOI21_X1 port map( B1 => n5926, B2 => n10226, A => n13788, ZN => 
                           n13783);
   U12327 : NAND3_X1 port map( A1 => n13789, A2 => n13790, A3 => n13791, ZN => 
                           n11904);
   U12328 : AOI221_X1 port map( B1 => n13792, B2 => n4863, C1 => n13793, C2 => 
                           MEM_IN(0), A => n13794, ZN => n13791);
   U12329 : OAI22_X1 port map( A1 => n10541, A2 => n251, B1 => n4867, B2 => 
                           n121, ZN => n13794);
   U12330 : NOR2_X1 port map( A1 => n5534, A2 => n13796, ZN => n5531);
   U12331 : INV_X1 port map( A => MEM_IN(0), ZN => n5534);
   U12332 : AOI22_X1 port map( A1 => n197, A2 => n4869, B1 => n150, B2 => n4871
                           , ZN => n13790);
   U12333 : NOR4_X1 port map( A1 => n13799, A2 => n13800, A3 => n13801, A4 => 
                           n13802, ZN => n13798);
   U12334 : OAI221_X1 port map( B1 => n11117, B2 => n316, C1 => n11053, C2 => 
                           n327, A => n13805, ZN => n13802);
   U12335 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_15_0_port, B1 => 
                           n13807, B2 => REGISTERS_11_0_port, C1 => n13808, C2 
                           => REGISTERS_39_0_port, ZN => n13805);
   U12336 : OAI221_X1 port map( B1 => n10829, B2 => n13809, C1 => n10957, C2 =>
                           n13810, A => n13811, ZN => n13801);
   U12337 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_0_port, B1 => 
                           n13813, B2 => REGISTERS_6_0_port, C1 => n347, C2 => 
                           REGISTERS_10_0_port, ZN => n13811);
   U12338 : OAI221_X1 port map( B1 => n10669, B2 => n13815, C1 => n10797, C2 =>
                           n303, A => n13817, ZN => n13800);
   U12339 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_0_port, B1 => 
                           n13819, B2 => REGISTERS_2_0_port, C1 => n358, C2 => 
                           REGISTERS_5_0_port, ZN => n13817);
   U12340 : OAI221_X1 port map( B1 => n10637, B2 => n13821, C1 => n11661, C2 =>
                           n304, A => n13823, ZN => n13799);
   U12341 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_0_port, B1 => 
                           n13825, B2 => REGISTERS_0_0_port, C1 => n13826, C2 
                           => REGISTERS_1_0_port, ZN => n13823);
   U12342 : NOR4_X1 port map( A1 => n13827, A2 => n13828, A3 => n13829, A4 => 
                           n13830, ZN => n13797);
   U12343 : OAI221_X1 port map( B1 => n11725, B2 => n371, C1 => n10989, C2 => 
                           n382, A => n13833_port, ZN => n13830);
   U12344 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_30_0_port, B1 => 
                           n404, B2 => REGISTERS_34_0_port, C1 => n415, C2 => 
                           REGISTERS_38_0_port, ZN => n13833_port);
   U12345 : OAI221_X1 port map( B1 => n11565, B2 => n426, C1 => n11693, C2 => 
                           n437, A => n13839_port, ZN => n13829);
   U12346 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_25_0_port, B1 => 
                           n459, B2 => REGISTERS_29_0_port, C1 => n470, C2 => 
                           REGISTERS_33_0_port, ZN => n13839_port);
   U12347 : OAI221_X1 port map( B1 => n11405, B2 => n481, C1 => n11533, C2 => 
                           n492, A => n13845_port, ZN => n13828);
   U12348 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_20_0_port, B1 => 
                           n514, B2 => REGISTERS_24_0_port, C1 => n525, C2 => 
                           REGISTERS_28_0_port, ZN => n13845_port);
   U12349 : OAI221_X1 port map( B1 => n11245, B2 => n536, C1 => n11373, C2 => 
                           n547, A => n13851_port, ZN => n13827);
   U12350 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_23_0_port, B1 => 
                           n569, B2 => REGISTERS_21_0_port, C1 => n580, C2 => 
                           REGISTERS_19_0_port, ZN => n13851_port);
   U12351 : NOR4_X1 port map( A1 => n13857_port, A2 => n13858_port, A3 => 
                           n13859_port, A4 => n13860_port, ZN => n13856_port);
   U12352 : OAI221_X1 port map( B1 => n11149, B2 => n316, C1 => n11085, C2 => 
                           n327, A => n13861_port, ZN => n13860_port);
   U12353 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_16_0_port, B1 => 
                           n119, B2 => REGISTERS_14_0_port, C1 => n13807, C2 =>
                           REGISTERS_12_0_port, ZN => n13861_port);
   U12354 : OAI221_X1 port map( B1 => n11117, B2 => n13863, C1 => n10861, C2 =>
                           n13809, A => n13864, ZN => n13859_port);
   U12355 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_0_port, B1 => 
                           n13865, B2 => REGISTERS_9_0_port, C1 => n13813, C2 
                           => REGISTERS_7_0_port, ZN => n13864);
   U12356 : OAI221_X1 port map( B1 => n10957, B2 => n13866, C1 => n10701, C2 =>
                           n13815, A => n13867, ZN => n13858_port);
   U12357 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_0_port, B1 => 
                           n13868, B2 => REGISTERS_36_0_port, C1 => n13819, C2 
                           => REGISTERS_3_0_port, ZN => n13867);
   U12358 : OAI221_X1 port map( B1 => n10797, B2 => n13869, C1 => n10669, C2 =>
                           n13821, A => n13870, ZN => n13857_port);
   U12359 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_0_port, B1 => 
                           n13871, B2 => REGISTERS_0_0_port, C1 => n13825, C2 
                           => REGISTERS_1_0_port, ZN => n13870);
   U12360 : NOR4_X1 port map( A1 => n13872, A2 => n13873, A3 => n13874, A4 => 
                           n13875, ZN => n13855_port);
   U12361 : OAI221_X1 port map( B1 => n11757, B2 => n371, C1 => n11021, C2 => 
                           n382, A => n13876, ZN => n13875);
   U12362 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_31_0_port, B1 => 
                           n404, B2 => REGISTERS_35_0_port, C1 => n415, C2 => 
                           REGISTERS_39_0_port, ZN => n13876);
   U12363 : OAI221_X1 port map( B1 => n11597, B2 => n426, C1 => n11725, C2 => 
                           n437, A => n13877, ZN => n13874);
   U12364 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_26_0_port, B1 => 
                           n459, B2 => REGISTERS_30_0_port, C1 => n470, C2 => 
                           REGISTERS_34_0_port, ZN => n13877);
   U12365 : OAI221_X1 port map( B1 => n11437, B2 => n481, C1 => n11565, C2 => 
                           n492, A => n13878, ZN => n13873);
   U12366 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_21_0_port, B1 => 
                           n514, B2 => REGISTERS_25_0_port, C1 => n525, C2 => 
                           REGISTERS_29_0_port, ZN => n13878);
   U12367 : OAI221_X1 port map( B1 => n11277, B2 => n536, C1 => n11405, C2 => 
                           n547, A => n13879, ZN => n13872);
   U12368 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_24_0_port, B1 => 
                           n569, B2 => REGISTERS_22_0_port, C1 => n580, C2 => 
                           REGISTERS_20_0_port, ZN => n13879);
   U12369 : AOI22_X1 port map( A1 => n13880, A2 => n4873, B1 => n13881, B2 => 
                           n4875, ZN => n13789);
   U12370 : NOR4_X1 port map( A1 => n13884, A2 => n13885, A3 => n13886, A4 => 
                           n13887, ZN => n13883);
   U12371 : OAI221_X1 port map( B1 => n11085, B2 => n316, C1 => n11021, C2 => 
                           n327, A => n13888, ZN => n13887);
   U12372 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_14_0_port, B1 => 
                           n13808, B2 => REGISTERS_38_0_port, C1 => n13889, C2 
                           => REGISTERS_39_0_port, ZN => n13888);
   U12373 : OAI221_X1 port map( B1 => n10925, B2 => n13810, C1 => n10861, C2 =>
                           n13890, A => n13891, ZN => n13886);
   U12374 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_0_port, B1 => 
                           n346, B2 => REGISTERS_9_0_port, C1 => n13812, C2 => 
                           REGISTERS_16_0_port, ZN => n13891);
   U12375 : OAI221_X1 port map( B1 => n10765, B2 => n303, C1 => n10701, C2 => 
                           n13893, A => n13894, ZN => n13885);
   U12376 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_0_port, B1 => 
                           n357, B2 => REGISTERS_4_0_port, C1 => n13818, C2 => 
                           REGISTERS_11_0_port, ZN => n13894);
   U12377 : OAI221_X1 port map( B1 => n11629, B2 => n304, C1 => n10573, C2 => 
                           n13896, A => n13897, ZN => n13884);
   U12378 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_0_port, B1 => 
                           n13826, B2 => REGISTERS_0_0_port, C1 => n13824, C2 
                           => REGISTERS_6_0_port, ZN => n13897);
   U12379 : NOR4_X1 port map( A1 => n13899, A2 => n13900, A3 => n13901, A4 => 
                           n13902, ZN => n13882);
   U12380 : OAI221_X1 port map( B1 => n11693, B2 => n371, C1 => n10957, C2 => 
                           n382, A => n13903, ZN => n13902);
   U12381 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_29_0_port, B1 => 
                           n404, B2 => REGISTERS_33_0_port, C1 => n415, C2 => 
                           REGISTERS_37_0_port, ZN => n13903);
   U12382 : OAI221_X1 port map( B1 => n11533, B2 => n426, C1 => n11661, C2 => 
                           n437, A => n13904, ZN => n13901);
   U12383 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_24_0_port, B1 => 
                           n459, B2 => REGISTERS_28_0_port, C1 => n470, C2 => 
                           REGISTERS_32_0_port, ZN => n13904);
   U12384 : OAI221_X1 port map( B1 => n11373, B2 => n481, C1 => n11501, C2 => 
                           n492, A => n13905, ZN => n13900);
   U12385 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_19_0_port, B1 => 
                           n514, B2 => REGISTERS_23_0_port, C1 => n525, C2 => 
                           REGISTERS_27_0_port, ZN => n13905);
   U12386 : OAI221_X1 port map( B1 => n11213, B2 => n536, C1 => n11341, C2 => 
                           n547, A => n13906, ZN => n13899);
   U12387 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_22_0_port, B1 => 
                           n569, B2 => REGISTERS_20_0_port, C1 => n580, C2 => 
                           REGISTERS_18_0_port, ZN => n13906);
   U12388 : NOR4_X1 port map( A1 => n13909, A2 => n13910, A3 => n13911, A4 => 
                           n13912, ZN => n13908);
   U12389 : OAI221_X1 port map( B1 => n11053, B2 => n316, C1 => n10989, C2 => 
                           n327, A => n13913, ZN => n13912);
   U12390 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_13_0_port, B1 => 
                           n13808, B2 => REGISTERS_37_0_port, C1 => n13889, C2 
                           => REGISTERS_38_0_port, ZN => n13913);
   U12391 : OAI221_X1 port map( B1 => n10893, B2 => n13810, C1 => n10829, C2 =>
                           n13890, A => n13914, ZN => n13911);
   U12392 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_0_port, B1 => 
                           n346, B2 => REGISTERS_8_0_port, C1 => n13812, C2 => 
                           REGISTERS_15_0_port, ZN => n13914);
   U12393 : OAI221_X1 port map( B1 => n10733, B2 => n303, C1 => n10669, C2 => 
                           n13893, A => n13915, ZN => n13910);
   U12394 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_0_port, B1 => 
                           n357, B2 => REGISTERS_3_0_port, C1 => n13818, C2 => 
                           REGISTERS_10_0_port, ZN => n13915);
   U12395 : OAI221_X1 port map( B1 => n11597, B2 => n304, C1 => n10541, C2 => 
                           n13896, A => n13916, ZN => n13909);
   U12396 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_0_port, B1 => 
                           n13917, B2 => REGISTERS_39_0_port, C1 => n13824, C2 
                           => REGISTERS_5_0_port, ZN => n13916);
   U12397 : NOR4_X1 port map( A1 => n13918, A2 => n13919, A3 => n13920, A4 => 
                           n13921, ZN => n13907);
   U12398 : OAI221_X1 port map( B1 => n11661, B2 => n371, C1 => n10925, C2 => 
                           n382, A => n13922, ZN => n13921);
   U12399 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_28_0_port, B1 => 
                           n404, B2 => REGISTERS_32_0_port, C1 => n415, C2 => 
                           REGISTERS_36_0_port, ZN => n13922);
   U12400 : OAI221_X1 port map( B1 => n11501, B2 => n426, C1 => n11629, C2 => 
                           n437, A => n13923, ZN => n13920);
   U12401 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_23_0_port, B1 => 
                           n459, B2 => REGISTERS_27_0_port, C1 => n470, C2 => 
                           REGISTERS_31_0_port, ZN => n13923);
   U12402 : OAI221_X1 port map( B1 => n11341, B2 => n481, C1 => n11469, C2 => 
                           n492, A => n13924, ZN => n13919);
   U12403 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_18_0_port, B1 => 
                           n514, B2 => REGISTERS_22_0_port, C1 => n525, C2 => 
                           REGISTERS_26_0_port, ZN => n13924);
   U12404 : OAI221_X1 port map( B1 => n11181, B2 => n536, C1 => n11309, C2 => 
                           n547, A => n13925, ZN => n13918);
   U12405 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_21_0_port, B1 => 
                           n569, B2 => REGISTERS_19_0_port, C1 => n580, C2 => 
                           REGISTERS_17_0_port, ZN => n13925);
   U12406 : NAND3_X1 port map( A1 => n13926, A2 => n13927, A3 => n13928, ZN => 
                           n11903);
   U12407 : AOI221_X1 port map( B1 => n13792, B2 => n4879, C1 => n13793, C2 => 
                           MEM_IN(1), A => n13929, ZN => n13928);
   U12408 : OAI22_X1 port map( A1 => n10538, A2 => n251, B1 => n4881, B2 => 
                           n121, ZN => n13929);
   U12409 : NOR2_X1 port map( A1 => n5543, A2 => n13796, ZN => n5541);
   U12410 : INV_X1 port map( A => MEM_IN(1), ZN => n5543);
   U12411 : AOI22_X1 port map( A1 => n197, A2 => n4882, B1 => n150, B2 => n4883
                           , ZN => n13927);
   U12412 : NOR4_X1 port map( A1 => n13932, A2 => n13933, A3 => n13934, A4 => 
                           n13935, ZN => n13931);
   U12413 : OAI221_X1 port map( B1 => n11116, B2 => n316, C1 => n11052, C2 => 
                           n327, A => n13936, ZN => n13935);
   U12414 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_15_1_port, B1 => 
                           n13807, B2 => REGISTERS_11_1_port, C1 => n13808, C2 
                           => REGISTERS_39_1_port, ZN => n13936);
   U12415 : OAI221_X1 port map( B1 => n10828, B2 => n13809, C1 => n10956, C2 =>
                           n13810, A => n13937, ZN => n13934);
   U12416 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_1_port, B1 => 
                           n13813, B2 => REGISTERS_6_1_port, C1 => n347, C2 => 
                           REGISTERS_10_1_port, ZN => n13937);
   U12417 : OAI221_X1 port map( B1 => n10668, B2 => n13815, C1 => n10796, C2 =>
                           n303, A => n13938, ZN => n13933);
   U12418 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_1_port, B1 => 
                           n13819, B2 => REGISTERS_2_1_port, C1 => n358, C2 => 
                           REGISTERS_5_1_port, ZN => n13938);
   U12419 : OAI221_X1 port map( B1 => n10636, B2 => n13821, C1 => n11660, C2 =>
                           n304, A => n13939, ZN => n13932);
   U12420 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_1_port, B1 => 
                           n13825, B2 => REGISTERS_0_1_port, C1 => n13826, C2 
                           => REGISTERS_1_1_port, ZN => n13939);
   U12421 : NOR4_X1 port map( A1 => n13940, A2 => n13941, A3 => n13942, A4 => 
                           n13943, ZN => n13930);
   U12422 : OAI221_X1 port map( B1 => n11724, B2 => n371, C1 => n10988, C2 => 
                           n382, A => n13944, ZN => n13943);
   U12423 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_30_1_port, B1 => 
                           n404, B2 => REGISTERS_34_1_port, C1 => n415, C2 => 
                           REGISTERS_38_1_port, ZN => n13944);
   U12424 : OAI221_X1 port map( B1 => n11564, B2 => n426, C1 => n11692, C2 => 
                           n437, A => n13945, ZN => n13942);
   U12425 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_25_1_port, B1 => 
                           n459, B2 => REGISTERS_29_1_port, C1 => n470, C2 => 
                           REGISTERS_33_1_port, ZN => n13945);
   U12426 : OAI221_X1 port map( B1 => n11404, B2 => n481, C1 => n11532, C2 => 
                           n492, A => n13946, ZN => n13941);
   U12427 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_20_1_port, B1 => 
                           n514, B2 => REGISTERS_24_1_port, C1 => n525, C2 => 
                           REGISTERS_28_1_port, ZN => n13946);
   U12428 : OAI221_X1 port map( B1 => n11244, B2 => n536, C1 => n11372, C2 => 
                           n547, A => n13947, ZN => n13940);
   U12429 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_23_1_port, B1 => 
                           n569, B2 => REGISTERS_21_1_port, C1 => n580, C2 => 
                           REGISTERS_19_1_port, ZN => n13947);
   U12430 : NOR4_X1 port map( A1 => n13950, A2 => n13951, A3 => n13952, A4 => 
                           n13953, ZN => n13949);
   U12431 : OAI221_X1 port map( B1 => n11148, B2 => n316, C1 => n11084, C2 => 
                           n327, A => n13954, ZN => n13953);
   U12432 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_16_1_port, B1 => 
                           n119, B2 => REGISTERS_14_1_port, C1 => n13807, C2 =>
                           REGISTERS_12_1_port, ZN => n13954);
   U12433 : OAI221_X1 port map( B1 => n11116, B2 => n13863, C1 => n10860, C2 =>
                           n13809, A => n13955, ZN => n13952);
   U12434 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_1_port, B1 => 
                           n13865, B2 => REGISTERS_9_1_port, C1 => n13813, C2 
                           => REGISTERS_7_1_port, ZN => n13955);
   U12435 : OAI221_X1 port map( B1 => n10956, B2 => n13866, C1 => n10700, C2 =>
                           n13815, A => n13956, ZN => n13951);
   U12436 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_1_port, B1 => 
                           n13868, B2 => REGISTERS_36_1_port, C1 => n13819, C2 
                           => REGISTERS_3_1_port, ZN => n13956);
   U12437 : OAI221_X1 port map( B1 => n10796, B2 => n13869, C1 => n10668, C2 =>
                           n13821, A => n13957, ZN => n13950);
   U12438 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_1_port, B1 => 
                           n13871, B2 => REGISTERS_0_1_port, C1 => n13825, C2 
                           => REGISTERS_1_1_port, ZN => n13957);
   U12439 : NOR4_X1 port map( A1 => n13958, A2 => n13959, A3 => n13960, A4 => 
                           n13961, ZN => n13948);
   U12440 : OAI221_X1 port map( B1 => n11756, B2 => n371, C1 => n11020, C2 => 
                           n382, A => n13962, ZN => n13961);
   U12441 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_31_1_port, B1 => 
                           n404, B2 => REGISTERS_35_1_port, C1 => n415, C2 => 
                           REGISTERS_39_1_port, ZN => n13962);
   U12442 : OAI221_X1 port map( B1 => n11596, B2 => n426, C1 => n11724, C2 => 
                           n437, A => n13963, ZN => n13960);
   U12443 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_26_1_port, B1 => 
                           n459, B2 => REGISTERS_30_1_port, C1 => n470, C2 => 
                           REGISTERS_34_1_port, ZN => n13963);
   U12444 : OAI221_X1 port map( B1 => n11436, B2 => n481, C1 => n11564, C2 => 
                           n492, A => n13964, ZN => n13959);
   U12445 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_21_1_port, B1 => 
                           n514, B2 => REGISTERS_25_1_port, C1 => n525, C2 => 
                           REGISTERS_29_1_port, ZN => n13964);
   U12446 : OAI221_X1 port map( B1 => n11276, B2 => n536, C1 => n11404, C2 => 
                           n547, A => n13965, ZN => n13958);
   U12447 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_24_1_port, B1 => 
                           n569, B2 => REGISTERS_22_1_port, C1 => n580, C2 => 
                           REGISTERS_20_1_port, ZN => n13965);
   U12448 : AOI22_X1 port map( A1 => n13880, A2 => n4884, B1 => n13881, B2 => 
                           n4885, ZN => n13926);
   U12449 : NOR4_X1 port map( A1 => n13968, A2 => n13969, A3 => n13970, A4 => 
                           n13971, ZN => n13967);
   U12450 : OAI221_X1 port map( B1 => n11084, B2 => n316, C1 => n11020, C2 => 
                           n327, A => n13972, ZN => n13971);
   U12451 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_14_1_port, B1 => 
                           n13808, B2 => REGISTERS_38_1_port, C1 => n13889, C2 
                           => REGISTERS_39_1_port, ZN => n13972);
   U12452 : OAI221_X1 port map( B1 => n10924, B2 => n13810, C1 => n10860, C2 =>
                           n13890, A => n13973, ZN => n13970);
   U12453 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_1_port, B1 => 
                           n345, B2 => REGISTERS_9_1_port, C1 => n13812, C2 => 
                           REGISTERS_16_1_port, ZN => n13973);
   U12454 : OAI221_X1 port map( B1 => n10764, B2 => n303, C1 => n10700, C2 => 
                           n13893, A => n13974, ZN => n13969);
   U12455 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_1_port, B1 => 
                           n356, B2 => REGISTERS_4_1_port, C1 => n13818, C2 => 
                           REGISTERS_11_1_port, ZN => n13974);
   U12456 : OAI221_X1 port map( B1 => n11628, B2 => n304, C1 => n10572, C2 => 
                           n13896, A => n13975, ZN => n13968);
   U12457 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_1_port, B1 => 
                           n13826, B2 => REGISTERS_0_1_port, C1 => n13824, C2 
                           => REGISTERS_6_1_port, ZN => n13975);
   U12458 : NOR4_X1 port map( A1 => n13976, A2 => n13977, A3 => n13978, A4 => 
                           n13979, ZN => n13966);
   U12459 : OAI221_X1 port map( B1 => n11692, B2 => n371, C1 => n10956, C2 => 
                           n382, A => n13980, ZN => n13979);
   U12460 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_29_1_port, B1 => 
                           n404, B2 => REGISTERS_33_1_port, C1 => n415, C2 => 
                           REGISTERS_37_1_port, ZN => n13980);
   U12461 : OAI221_X1 port map( B1 => n11532, B2 => n426, C1 => n11660, C2 => 
                           n437, A => n13981, ZN => n13978);
   U12462 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_24_1_port, B1 => 
                           n459, B2 => REGISTERS_28_1_port, C1 => n470, C2 => 
                           REGISTERS_32_1_port, ZN => n13981);
   U12463 : OAI221_X1 port map( B1 => n11372, B2 => n481, C1 => n11500, C2 => 
                           n492, A => n13982, ZN => n13977);
   U12464 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_19_1_port, B1 => 
                           n514, B2 => REGISTERS_23_1_port, C1 => n525, C2 => 
                           REGISTERS_27_1_port, ZN => n13982);
   U12465 : OAI221_X1 port map( B1 => n11212, B2 => n536, C1 => n11340, C2 => 
                           n547, A => n13983, ZN => n13976);
   U12466 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_22_1_port, B1 => 
                           n569, B2 => REGISTERS_20_1_port, C1 => n580, C2 => 
                           REGISTERS_18_1_port, ZN => n13983);
   U12467 : NOR4_X1 port map( A1 => n13986, A2 => n13987, A3 => n13988, A4 => 
                           n13989, ZN => n13985);
   U12468 : OAI221_X1 port map( B1 => n11052, B2 => n316, C1 => n10988, C2 => 
                           n327, A => n13990, ZN => n13989);
   U12469 : AOI222_X1 port map( A1 => n338, A2 => REGISTERS_13_1_port, B1 => 
                           n13808, B2 => REGISTERS_37_1_port, C1 => n13889, C2 
                           => REGISTERS_38_1_port, ZN => n13990);
   U12470 : OAI221_X1 port map( B1 => n10892, B2 => n13810, C1 => n10828, C2 =>
                           n13890, A => n13991, ZN => n13988);
   U12471 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_1_port, B1 => 
                           n345, B2 => REGISTERS_8_1_port, C1 => n13812, C2 => 
                           REGISTERS_15_1_port, ZN => n13991);
   U12472 : OAI221_X1 port map( B1 => n10732, B2 => n303, C1 => n10668, C2 => 
                           n13893, A => n13992, ZN => n13987);
   U12473 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_1_port, B1 => 
                           n356, B2 => REGISTERS_3_1_port, C1 => n13818, C2 => 
                           REGISTERS_10_1_port, ZN => n13992);
   U12474 : OAI221_X1 port map( B1 => n11596, B2 => n304, C1 => n10538, C2 => 
                           n13896, A => n13993, ZN => n13986);
   U12475 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_1_port, B1 => 
                           n13917, B2 => REGISTERS_39_1_port, C1 => n13824, C2 
                           => REGISTERS_5_1_port, ZN => n13993);
   U12476 : NOR4_X1 port map( A1 => n13994, A2 => n13995, A3 => n13996, A4 => 
                           n13997, ZN => n13984);
   U12477 : OAI221_X1 port map( B1 => n11660, B2 => n371, C1 => n10924, C2 => 
                           n382, A => n13998, ZN => n13997);
   U12478 : AOI222_X1 port map( A1 => n393, A2 => REGISTERS_28_1_port, B1 => 
                           n404, B2 => REGISTERS_32_1_port, C1 => n415, C2 => 
                           REGISTERS_36_1_port, ZN => n13998);
   U12479 : OAI221_X1 port map( B1 => n11500, B2 => n426, C1 => n11628, C2 => 
                           n437, A => n13999, ZN => n13996);
   U12480 : AOI222_X1 port map( A1 => n448, A2 => REGISTERS_23_1_port, B1 => 
                           n459, B2 => REGISTERS_27_1_port, C1 => n470, C2 => 
                           REGISTERS_31_1_port, ZN => n13999);
   U12481 : OAI221_X1 port map( B1 => n11340, B2 => n481, C1 => n11468, C2 => 
                           n492, A => n14000, ZN => n13995);
   U12482 : AOI222_X1 port map( A1 => n503, A2 => REGISTERS_18_1_port, B1 => 
                           n514, B2 => REGISTERS_22_1_port, C1 => n525, C2 => 
                           REGISTERS_26_1_port, ZN => n14000);
   U12483 : OAI221_X1 port map( B1 => n11180, B2 => n536, C1 => n11308, C2 => 
                           n547, A => n14001, ZN => n13994);
   U12484 : AOI222_X1 port map( A1 => n558, A2 => REGISTERS_21_1_port, B1 => 
                           n569, B2 => REGISTERS_19_1_port, C1 => n580, C2 => 
                           REGISTERS_17_1_port, ZN => n14001);
   U12485 : NAND3_X1 port map( A1 => n14002, A2 => n14003, A3 => n14004, ZN => 
                           n11902);
   U12486 : AOI221_X1 port map( B1 => n13792, B2 => n4889, C1 => n13793, C2 => 
                           MEM_IN(2), A => n14005, ZN => n14004);
   U12487 : OAI22_X1 port map( A1 => n10535, A2 => n251, B1 => n4891, B2 => 
                           n121, ZN => n14005);
   U12488 : NOR2_X1 port map( A1 => n5550, A2 => n13796, ZN => n5548);
   U12489 : INV_X1 port map( A => MEM_IN(2), ZN => n5550);
   U12490 : AOI22_X1 port map( A1 => n197, A2 => n4892, B1 => n150, B2 => n4893
                           , ZN => n14003);
   U12491 : NOR4_X1 port map( A1 => n14008, A2 => n14009, A3 => n14010, A4 => 
                           n14011, ZN => n14007);
   U12492 : OAI221_X1 port map( B1 => n11115, B2 => n315, C1 => n11051, C2 => 
                           n326, A => n14012, ZN => n14011);
   U12493 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_15_2_port, B1 => 
                           n13807, B2 => REGISTERS_11_2_port, C1 => n13808, C2 
                           => REGISTERS_39_2_port, ZN => n14012);
   U12494 : OAI221_X1 port map( B1 => n10827, B2 => n13809, C1 => n10955, C2 =>
                           n13810, A => n14013, ZN => n14010);
   U12495 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_2_port, B1 => 
                           n13813, B2 => REGISTERS_6_2_port, C1 => n347, C2 => 
                           REGISTERS_10_2_port, ZN => n14013);
   U12496 : OAI221_X1 port map( B1 => n10667, B2 => n13815, C1 => n10795, C2 =>
                           n303, A => n14014, ZN => n14009);
   U12497 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_2_port, B1 => 
                           n13819, B2 => REGISTERS_2_2_port, C1 => n358, C2 => 
                           REGISTERS_5_2_port, ZN => n14014);
   U12498 : OAI221_X1 port map( B1 => n10635, B2 => n13821, C1 => n11659, C2 =>
                           n304, A => n14015, ZN => n14008);
   U12499 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_2_port, B1 => 
                           n13825, B2 => REGISTERS_0_2_port, C1 => n13826, C2 
                           => REGISTERS_1_2_port, ZN => n14015);
   U12500 : NOR4_X1 port map( A1 => n14016, A2 => n14017, A3 => n14018, A4 => 
                           n14019, ZN => n14006);
   U12501 : OAI221_X1 port map( B1 => n11723, B2 => n370, C1 => n10987, C2 => 
                           n382, A => n14020, ZN => n14019);
   U12502 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_30_2_port, B1 => 
                           n403, B2 => REGISTERS_34_2_port, C1 => n414, C2 => 
                           REGISTERS_38_2_port, ZN => n14020);
   U12503 : OAI221_X1 port map( B1 => n11563, B2 => n425, C1 => n11691, C2 => 
                           n436, A => n14021, ZN => n14018);
   U12504 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_25_2_port, B1 => 
                           n458, B2 => REGISTERS_29_2_port, C1 => n469, C2 => 
                           REGISTERS_33_2_port, ZN => n14021);
   U12505 : OAI221_X1 port map( B1 => n11403, B2 => n480, C1 => n11531, C2 => 
                           n491, A => n14022, ZN => n14017);
   U12506 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_20_2_port, B1 => 
                           n513, B2 => REGISTERS_24_2_port, C1 => n524, C2 => 
                           REGISTERS_28_2_port, ZN => n14022);
   U12507 : OAI221_X1 port map( B1 => n11243, B2 => n535, C1 => n11371, C2 => 
                           n546, A => n14023, ZN => n14016);
   U12508 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_23_2_port, B1 => 
                           n568, B2 => REGISTERS_21_2_port, C1 => n579, C2 => 
                           REGISTERS_19_2_port, ZN => n14023);
   U12509 : NOR4_X1 port map( A1 => n14026, A2 => n14027, A3 => n14028, A4 => 
                           n14029, ZN => n14025);
   U12510 : OAI221_X1 port map( B1 => n11147, B2 => n315, C1 => n11083, C2 => 
                           n326, A => n14030, ZN => n14029);
   U12511 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_16_2_port, B1 => 
                           n119, B2 => REGISTERS_14_2_port, C1 => n13807, C2 =>
                           REGISTERS_12_2_port, ZN => n14030);
   U12512 : OAI221_X1 port map( B1 => n11115, B2 => n13863, C1 => n10859, C2 =>
                           n13809, A => n14031, ZN => n14028);
   U12513 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_2_port, B1 => 
                           n13865, B2 => REGISTERS_9_2_port, C1 => n13813, C2 
                           => REGISTERS_7_2_port, ZN => n14031);
   U12514 : OAI221_X1 port map( B1 => n10955, B2 => n13866, C1 => n10699, C2 =>
                           n13815, A => n14032, ZN => n14027);
   U12515 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_2_port, B1 => 
                           n13868, B2 => REGISTERS_36_2_port, C1 => n13819, C2 
                           => REGISTERS_3_2_port, ZN => n14032);
   U12516 : OAI221_X1 port map( B1 => n10795, B2 => n13869, C1 => n10667, C2 =>
                           n13821, A => n14033, ZN => n14026);
   U12517 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_2_port, B1 => 
                           n13871, B2 => REGISTERS_0_2_port, C1 => n13825, C2 
                           => REGISTERS_1_2_port, ZN => n14033);
   U12518 : NOR4_X1 port map( A1 => n14034, A2 => n14035, A3 => n14036, A4 => 
                           n14037, ZN => n14024);
   U12519 : OAI221_X1 port map( B1 => n11755, B2 => n370, C1 => n11019, C2 => 
                           n381, A => n14038, ZN => n14037);
   U12520 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_31_2_port, B1 => 
                           n403, B2 => REGISTERS_35_2_port, C1 => n414, C2 => 
                           REGISTERS_39_2_port, ZN => n14038);
   U12521 : OAI221_X1 port map( B1 => n11595, B2 => n425, C1 => n11723, C2 => 
                           n436, A => n14039, ZN => n14036);
   U12522 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_26_2_port, B1 => 
                           n458, B2 => REGISTERS_30_2_port, C1 => n469, C2 => 
                           REGISTERS_34_2_port, ZN => n14039);
   U12523 : OAI221_X1 port map( B1 => n11435, B2 => n480, C1 => n11563, C2 => 
                           n491, A => n14040, ZN => n14035);
   U12524 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_21_2_port, B1 => 
                           n513, B2 => REGISTERS_25_2_port, C1 => n524, C2 => 
                           REGISTERS_29_2_port, ZN => n14040);
   U12525 : OAI221_X1 port map( B1 => n11275, B2 => n535, C1 => n11403, C2 => 
                           n546, A => n14041, ZN => n14034);
   U12526 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_24_2_port, B1 => 
                           n568, B2 => REGISTERS_22_2_port, C1 => n579, C2 => 
                           REGISTERS_20_2_port, ZN => n14041);
   U12527 : AOI22_X1 port map( A1 => n13880, A2 => n4894, B1 => n13881, B2 => 
                           n4895, ZN => n14002);
   U12528 : NOR4_X1 port map( A1 => n14044, A2 => n14045, A3 => n14046, A4 => 
                           n14047, ZN => n14043);
   U12529 : OAI221_X1 port map( B1 => n11083, B2 => n315, C1 => n11019, C2 => 
                           n326, A => n14048, ZN => n14047);
   U12530 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_14_2_port, B1 => 
                           n13808, B2 => REGISTERS_38_2_port, C1 => n13889, C2 
                           => REGISTERS_39_2_port, ZN => n14048);
   U12531 : OAI221_X1 port map( B1 => n10923, B2 => n13810, C1 => n10859, C2 =>
                           n13890, A => n14049, ZN => n14046);
   U12532 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_2_port, B1 => 
                           n345, B2 => REGISTERS_9_2_port, C1 => n13812, C2 => 
                           REGISTERS_16_2_port, ZN => n14049);
   U12533 : OAI221_X1 port map( B1 => n10763, B2 => n303, C1 => n10699, C2 => 
                           n13893, A => n14050, ZN => n14045);
   U12534 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_2_port, B1 => 
                           n356, B2 => REGISTERS_4_2_port, C1 => n13818, C2 => 
                           REGISTERS_11_2_port, ZN => n14050);
   U12535 : OAI221_X1 port map( B1 => n11627, B2 => n304, C1 => n10571, C2 => 
                           n13896, A => n14051, ZN => n14044);
   U12536 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_2_port, B1 => 
                           n13826, B2 => REGISTERS_0_2_port, C1 => n13824, C2 
                           => REGISTERS_6_2_port, ZN => n14051);
   U12537 : NOR4_X1 port map( A1 => n14052, A2 => n14053, A3 => n14054, A4 => 
                           n14055, ZN => n14042);
   U12538 : OAI221_X1 port map( B1 => n11691, B2 => n370, C1 => n10955, C2 => 
                           n381, A => n14056, ZN => n14055);
   U12539 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_29_2_port, B1 => 
                           n403, B2 => REGISTERS_33_2_port, C1 => n414, C2 => 
                           REGISTERS_37_2_port, ZN => n14056);
   U12540 : OAI221_X1 port map( B1 => n11531, B2 => n425, C1 => n11659, C2 => 
                           n436, A => n14057, ZN => n14054);
   U12541 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_24_2_port, B1 => 
                           n458, B2 => REGISTERS_28_2_port, C1 => n469, C2 => 
                           REGISTERS_32_2_port, ZN => n14057);
   U12542 : OAI221_X1 port map( B1 => n11371, B2 => n480, C1 => n11499, C2 => 
                           n491, A => n14058, ZN => n14053);
   U12543 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_19_2_port, B1 => 
                           n513, B2 => REGISTERS_23_2_port, C1 => n524, C2 => 
                           REGISTERS_27_2_port, ZN => n14058);
   U12544 : OAI221_X1 port map( B1 => n11211, B2 => n535, C1 => n11339, C2 => 
                           n546, A => n14059, ZN => n14052);
   U12545 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_22_2_port, B1 => 
                           n568, B2 => REGISTERS_20_2_port, C1 => n579, C2 => 
                           REGISTERS_18_2_port, ZN => n14059);
   U12546 : NOR4_X1 port map( A1 => n14062, A2 => n14063, A3 => n14064, A4 => 
                           n14065, ZN => n14061);
   U12547 : OAI221_X1 port map( B1 => n11051, B2 => n315, C1 => n10987, C2 => 
                           n326, A => n14066, ZN => n14065);
   U12548 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_13_2_port, B1 => 
                           n13808, B2 => REGISTERS_37_2_port, C1 => n13889, C2 
                           => REGISTERS_38_2_port, ZN => n14066);
   U12549 : OAI221_X1 port map( B1 => n10891, B2 => n13810, C1 => n10827, C2 =>
                           n13890, A => n14067, ZN => n14064);
   U12550 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_2_port, B1 => 
                           n344, B2 => REGISTERS_8_2_port, C1 => n13812, C2 => 
                           REGISTERS_15_2_port, ZN => n14067);
   U12551 : OAI221_X1 port map( B1 => n10731, B2 => n303, C1 => n10667, C2 => 
                           n13893, A => n14068, ZN => n14063);
   U12552 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_2_port, B1 => 
                           n355, B2 => REGISTERS_3_2_port, C1 => n13818, C2 => 
                           REGISTERS_10_2_port, ZN => n14068);
   U12553 : OAI221_X1 port map( B1 => n11595, B2 => n304, C1 => n10535, C2 => 
                           n13896, A => n14069, ZN => n14062);
   U12554 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_2_port, B1 => 
                           n13917, B2 => REGISTERS_39_2_port, C1 => n13824, C2 
                           => REGISTERS_5_2_port, ZN => n14069);
   U12555 : NOR4_X1 port map( A1 => n14070, A2 => n14071, A3 => n14072, A4 => 
                           n14073, ZN => n14060);
   U12556 : OAI221_X1 port map( B1 => n11659, B2 => n370, C1 => n10923, C2 => 
                           n381, A => n14074, ZN => n14073);
   U12557 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_28_2_port, B1 => 
                           n403, B2 => REGISTERS_32_2_port, C1 => n414, C2 => 
                           REGISTERS_36_2_port, ZN => n14074);
   U12558 : OAI221_X1 port map( B1 => n11499, B2 => n425, C1 => n11627, C2 => 
                           n436, A => n14075, ZN => n14072);
   U12559 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_23_2_port, B1 => 
                           n458, B2 => REGISTERS_27_2_port, C1 => n469, C2 => 
                           REGISTERS_31_2_port, ZN => n14075);
   U12560 : OAI221_X1 port map( B1 => n11339, B2 => n480, C1 => n11467, C2 => 
                           n491, A => n14076, ZN => n14071);
   U12561 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_18_2_port, B1 => 
                           n513, B2 => REGISTERS_22_2_port, C1 => n524, C2 => 
                           REGISTERS_26_2_port, ZN => n14076);
   U12562 : OAI221_X1 port map( B1 => n11179, B2 => n535, C1 => n11307, C2 => 
                           n546, A => n14077, ZN => n14070);
   U12563 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_21_2_port, B1 => 
                           n568, B2 => REGISTERS_19_2_port, C1 => n579, C2 => 
                           REGISTERS_17_2_port, ZN => n14077);
   U12564 : NAND3_X1 port map( A1 => n14078, A2 => n14079, A3 => n14080, ZN => 
                           n11901);
   U12565 : AOI221_X1 port map( B1 => n13792, B2 => n4899, C1 => n13793, C2 => 
                           MEM_IN(3), A => n14081, ZN => n14080);
   U12566 : OAI22_X1 port map( A1 => n10532, A2 => n251, B1 => n4901, B2 => 
                           n121, ZN => n14081);
   U12567 : NOR2_X1 port map( A1 => n5557, A2 => n13796, ZN => n5555);
   U12568 : INV_X1 port map( A => MEM_IN(3), ZN => n5557);
   U12569 : AOI22_X1 port map( A1 => n197, A2 => n4902, B1 => n150, B2 => n4903
                           , ZN => n14079);
   U12570 : NOR4_X1 port map( A1 => n14084, A2 => n14085, A3 => n14086, A4 => 
                           n14087, ZN => n14083);
   U12571 : OAI221_X1 port map( B1 => n11114, B2 => n315, C1 => n11050, C2 => 
                           n326, A => n14088, ZN => n14087);
   U12572 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_15_3_port, B1 => 
                           n13807, B2 => REGISTERS_11_3_port, C1 => n13808, C2 
                           => REGISTERS_39_3_port, ZN => n14088);
   U12573 : OAI221_X1 port map( B1 => n10826, B2 => n13809, C1 => n10954, C2 =>
                           n13810, A => n14089, ZN => n14086);
   U12574 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_3_port, B1 => 
                           n13813, B2 => REGISTERS_6_3_port, C1 => n347, C2 => 
                           REGISTERS_10_3_port, ZN => n14089);
   U12575 : OAI221_X1 port map( B1 => n10666, B2 => n13815, C1 => n10794, C2 =>
                           n303, A => n14090, ZN => n14085);
   U12576 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_3_port, B1 => 
                           n13819, B2 => REGISTERS_2_3_port, C1 => n358, C2 => 
                           REGISTERS_5_3_port, ZN => n14090);
   U12577 : OAI221_X1 port map( B1 => n10634, B2 => n13821, C1 => n11658, C2 =>
                           n304, A => n14091, ZN => n14084);
   U12578 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_3_port, B1 => 
                           n13825, B2 => REGISTERS_0_3_port, C1 => n13826, C2 
                           => REGISTERS_1_3_port, ZN => n14091);
   U12579 : NOR4_X1 port map( A1 => n14092, A2 => n14093, A3 => n14094, A4 => 
                           n14095, ZN => n14082);
   U12580 : OAI221_X1 port map( B1 => n11722, B2 => n370, C1 => n10986, C2 => 
                           n381, A => n14096, ZN => n14095);
   U12581 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_30_3_port, B1 => 
                           n403, B2 => REGISTERS_34_3_port, C1 => n414, C2 => 
                           REGISTERS_38_3_port, ZN => n14096);
   U12582 : OAI221_X1 port map( B1 => n11562, B2 => n425, C1 => n11690, C2 => 
                           n436, A => n14097, ZN => n14094);
   U12583 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_25_3_port, B1 => 
                           n458, B2 => REGISTERS_29_3_port, C1 => n469, C2 => 
                           REGISTERS_33_3_port, ZN => n14097);
   U12584 : OAI221_X1 port map( B1 => n11402, B2 => n480, C1 => n11530, C2 => 
                           n491, A => n14098, ZN => n14093);
   U12585 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_20_3_port, B1 => 
                           n513, B2 => REGISTERS_24_3_port, C1 => n524, C2 => 
                           REGISTERS_28_3_port, ZN => n14098);
   U12586 : OAI221_X1 port map( B1 => n11242, B2 => n535, C1 => n11370, C2 => 
                           n546, A => n14099, ZN => n14092);
   U12587 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_23_3_port, B1 => 
                           n568, B2 => REGISTERS_21_3_port, C1 => n579, C2 => 
                           REGISTERS_19_3_port, ZN => n14099);
   U12588 : NOR4_X1 port map( A1 => n14102, A2 => n14103, A3 => n14104, A4 => 
                           n14105, ZN => n14101);
   U12589 : OAI221_X1 port map( B1 => n11146, B2 => n315, C1 => n11082, C2 => 
                           n326, A => n14106, ZN => n14105);
   U12590 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_16_3_port, B1 => 
                           n119, B2 => REGISTERS_14_3_port, C1 => n13807, C2 =>
                           REGISTERS_12_3_port, ZN => n14106);
   U12591 : OAI221_X1 port map( B1 => n11114, B2 => n13863, C1 => n10858, C2 =>
                           n13809, A => n14107, ZN => n14104);
   U12592 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_3_port, B1 => 
                           n13865, B2 => REGISTERS_9_3_port, C1 => n13813, C2 
                           => REGISTERS_7_3_port, ZN => n14107);
   U12593 : OAI221_X1 port map( B1 => n10954, B2 => n13866, C1 => n10698, C2 =>
                           n13815, A => n14108, ZN => n14103);
   U12594 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_3_port, B1 => 
                           n13868, B2 => REGISTERS_36_3_port, C1 => n13819, C2 
                           => REGISTERS_3_3_port, ZN => n14108);
   U12595 : OAI221_X1 port map( B1 => n10794, B2 => n13869, C1 => n10666, C2 =>
                           n13821, A => n14109, ZN => n14102);
   U12596 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_3_port, B1 => 
                           n13871, B2 => REGISTERS_0_3_port, C1 => n13825, C2 
                           => REGISTERS_1_3_port, ZN => n14109);
   U12597 : NOR4_X1 port map( A1 => n14110, A2 => n14111, A3 => n14112, A4 => 
                           n14113, ZN => n14100);
   U12598 : OAI221_X1 port map( B1 => n11754, B2 => n370, C1 => n11018, C2 => 
                           n381, A => n14114, ZN => n14113);
   U12599 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_31_3_port, B1 => 
                           n403, B2 => REGISTERS_35_3_port, C1 => n414, C2 => 
                           REGISTERS_39_3_port, ZN => n14114);
   U12600 : OAI221_X1 port map( B1 => n11594, B2 => n425, C1 => n11722, C2 => 
                           n436, A => n14115, ZN => n14112);
   U12601 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_26_3_port, B1 => 
                           n458, B2 => REGISTERS_30_3_port, C1 => n469, C2 => 
                           REGISTERS_34_3_port, ZN => n14115);
   U12602 : OAI221_X1 port map( B1 => n11434, B2 => n480, C1 => n11562, C2 => 
                           n491, A => n14116, ZN => n14111);
   U12603 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_21_3_port, B1 => 
                           n513, B2 => REGISTERS_25_3_port, C1 => n524, C2 => 
                           REGISTERS_29_3_port, ZN => n14116);
   U12604 : OAI221_X1 port map( B1 => n11274, B2 => n535, C1 => n11402, C2 => 
                           n546, A => n14117, ZN => n14110);
   U12605 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_24_3_port, B1 => 
                           n568, B2 => REGISTERS_22_3_port, C1 => n579, C2 => 
                           REGISTERS_20_3_port, ZN => n14117);
   U12606 : AOI22_X1 port map( A1 => n13880, A2 => n4904, B1 => n13881, B2 => 
                           n4905, ZN => n14078);
   U12607 : NOR4_X1 port map( A1 => n14120, A2 => n14121, A3 => n14122, A4 => 
                           n14123, ZN => n14119);
   U12608 : OAI221_X1 port map( B1 => n11082, B2 => n315, C1 => n11018, C2 => 
                           n326, A => n14124, ZN => n14123);
   U12609 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_14_3_port, B1 => 
                           n13808, B2 => REGISTERS_38_3_port, C1 => n13889, C2 
                           => REGISTERS_39_3_port, ZN => n14124);
   U12610 : OAI221_X1 port map( B1 => n10922, B2 => n13810, C1 => n10858, C2 =>
                           n13890, A => n14125, ZN => n14122);
   U12611 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_3_port, B1 => 
                           n344, B2 => REGISTERS_9_3_port, C1 => n13812, C2 => 
                           REGISTERS_16_3_port, ZN => n14125);
   U12612 : OAI221_X1 port map( B1 => n10762, B2 => n303, C1 => n10698, C2 => 
                           n13893, A => n14126, ZN => n14121);
   U12613 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_3_port, B1 => 
                           n355, B2 => REGISTERS_4_3_port, C1 => n13818, C2 => 
                           REGISTERS_11_3_port, ZN => n14126);
   U12614 : OAI221_X1 port map( B1 => n11626, B2 => n304, C1 => n10570, C2 => 
                           n13896, A => n14127, ZN => n14120);
   U12615 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_3_port, B1 => 
                           n13826, B2 => REGISTERS_0_3_port, C1 => n13824, C2 
                           => REGISTERS_6_3_port, ZN => n14127);
   U12616 : NOR4_X1 port map( A1 => n14128, A2 => n14129, A3 => n14130, A4 => 
                           n14131, ZN => n14118);
   U12617 : OAI221_X1 port map( B1 => n11690, B2 => n370, C1 => n10954, C2 => 
                           n381, A => n14132, ZN => n14131);
   U12618 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_29_3_port, B1 => 
                           n403, B2 => REGISTERS_33_3_port, C1 => n414, C2 => 
                           REGISTERS_37_3_port, ZN => n14132);
   U12619 : OAI221_X1 port map( B1 => n11530, B2 => n425, C1 => n11658, C2 => 
                           n436, A => n14133, ZN => n14130);
   U12620 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_24_3_port, B1 => 
                           n458, B2 => REGISTERS_28_3_port, C1 => n469, C2 => 
                           REGISTERS_32_3_port, ZN => n14133);
   U12621 : OAI221_X1 port map( B1 => n11370, B2 => n480, C1 => n11498, C2 => 
                           n491, A => n14134, ZN => n14129);
   U12622 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_19_3_port, B1 => 
                           n513, B2 => REGISTERS_23_3_port, C1 => n524, C2 => 
                           REGISTERS_27_3_port, ZN => n14134);
   U12623 : OAI221_X1 port map( B1 => n11210, B2 => n535, C1 => n11338, C2 => 
                           n546, A => n14135, ZN => n14128);
   U12624 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_22_3_port, B1 => 
                           n568, B2 => REGISTERS_20_3_port, C1 => n579, C2 => 
                           REGISTERS_18_3_port, ZN => n14135);
   U12625 : NOR4_X1 port map( A1 => n14138, A2 => n14139, A3 => n14140, A4 => 
                           n14141, ZN => n14137);
   U12626 : OAI221_X1 port map( B1 => n11050, B2 => n315, C1 => n10986, C2 => 
                           n326, A => n14142, ZN => n14141);
   U12627 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_13_3_port, B1 => 
                           n13808, B2 => REGISTERS_37_3_port, C1 => n13889, C2 
                           => REGISTERS_38_3_port, ZN => n14142);
   U12628 : OAI221_X1 port map( B1 => n10890, B2 => n13810, C1 => n10826, C2 =>
                           n13890, A => n14143, ZN => n14140);
   U12629 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_3_port, B1 => 
                           n343, B2 => REGISTERS_8_3_port, C1 => n13812, C2 => 
                           REGISTERS_15_3_port, ZN => n14143);
   U12630 : OAI221_X1 port map( B1 => n10730, B2 => n303, C1 => n10666, C2 => 
                           n13893, A => n14144, ZN => n14139);
   U12631 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_3_port, B1 => 
                           n354, B2 => REGISTERS_3_3_port, C1 => n13818, C2 => 
                           REGISTERS_10_3_port, ZN => n14144);
   U12632 : OAI221_X1 port map( B1 => n11594, B2 => n304, C1 => n10532, C2 => 
                           n13896, A => n14145, ZN => n14138);
   U12633 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_3_port, B1 => 
                           n13917, B2 => REGISTERS_39_3_port, C1 => n13824, C2 
                           => REGISTERS_5_3_port, ZN => n14145);
   U12634 : NOR4_X1 port map( A1 => n14146, A2 => n14147, A3 => n14148, A4 => 
                           n14149, ZN => n14136);
   U12635 : OAI221_X1 port map( B1 => n11658, B2 => n370, C1 => n10922, C2 => 
                           n381, A => n14150, ZN => n14149);
   U12636 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_28_3_port, B1 => 
                           n403, B2 => REGISTERS_32_3_port, C1 => n414, C2 => 
                           REGISTERS_36_3_port, ZN => n14150);
   U12637 : OAI221_X1 port map( B1 => n11498, B2 => n425, C1 => n11626, C2 => 
                           n436, A => n14151, ZN => n14148);
   U12638 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_23_3_port, B1 => 
                           n458, B2 => REGISTERS_27_3_port, C1 => n469, C2 => 
                           REGISTERS_31_3_port, ZN => n14151);
   U12639 : OAI221_X1 port map( B1 => n11338, B2 => n480, C1 => n11466, C2 => 
                           n491, A => n14152, ZN => n14147);
   U12640 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_18_3_port, B1 => 
                           n513, B2 => REGISTERS_22_3_port, C1 => n524, C2 => 
                           REGISTERS_26_3_port, ZN => n14152);
   U12641 : OAI221_X1 port map( B1 => n11178, B2 => n535, C1 => n11306, C2 => 
                           n546, A => n14153, ZN => n14146);
   U12642 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_21_3_port, B1 => 
                           n568, B2 => REGISTERS_19_3_port, C1 => n579, C2 => 
                           REGISTERS_17_3_port, ZN => n14153);
   U12643 : NAND3_X1 port map( A1 => n14154, A2 => n14155, A3 => n14156, ZN => 
                           n11900);
   U12644 : AOI221_X1 port map( B1 => n13792, B2 => n4909, C1 => n13793, C2 => 
                           MEM_IN(4), A => n14157, ZN => n14156);
   U12645 : OAI22_X1 port map( A1 => n10529, A2 => n251, B1 => n4911, B2 => 
                           n121, ZN => n14157);
   U12646 : NOR2_X1 port map( A1 => n5564, A2 => n13796, ZN => n5562);
   U12647 : INV_X1 port map( A => MEM_IN(4), ZN => n5564);
   U12648 : AOI22_X1 port map( A1 => n197, A2 => n4912, B1 => n150, B2 => n4913
                           , ZN => n14155);
   U12649 : NOR4_X1 port map( A1 => n14160, A2 => n14161, A3 => n14162, A4 => 
                           n14163, ZN => n14159);
   U12650 : OAI221_X1 port map( B1 => n11113, B2 => n315, C1 => n11049, C2 => 
                           n326, A => n14164, ZN => n14163);
   U12651 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_15_4_port, B1 => 
                           n13807, B2 => REGISTERS_11_4_port, C1 => n13808, C2 
                           => REGISTERS_39_4_port, ZN => n14164);
   U12652 : OAI221_X1 port map( B1 => n10825, B2 => n13809, C1 => n10953, C2 =>
                           n13810, A => n14165, ZN => n14162);
   U12653 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_4_port, B1 => 
                           n13813, B2 => REGISTERS_6_4_port, C1 => n347, C2 => 
                           REGISTERS_10_4_port, ZN => n14165);
   U12654 : OAI221_X1 port map( B1 => n10665, B2 => n13815, C1 => n10793, C2 =>
                           n303, A => n14166, ZN => n14161);
   U12655 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_4_port, B1 => 
                           n13819, B2 => REGISTERS_2_4_port, C1 => n358, C2 => 
                           REGISTERS_5_4_port, ZN => n14166);
   U12656 : OAI221_X1 port map( B1 => n10633, B2 => n13821, C1 => n11657, C2 =>
                           n304, A => n14167, ZN => n14160);
   U12657 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_4_port, B1 => 
                           n13825, B2 => REGISTERS_0_4_port, C1 => n13826, C2 
                           => REGISTERS_1_4_port, ZN => n14167);
   U12658 : NOR4_X1 port map( A1 => n14168, A2 => n14169, A3 => n14170, A4 => 
                           n14171, ZN => n14158);
   U12659 : OAI221_X1 port map( B1 => n11721, B2 => n370, C1 => n10985, C2 => 
                           n381, A => n14172, ZN => n14171);
   U12660 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_30_4_port, B1 => 
                           n403, B2 => REGISTERS_34_4_port, C1 => n414, C2 => 
                           REGISTERS_38_4_port, ZN => n14172);
   U12661 : OAI221_X1 port map( B1 => n11561, B2 => n425, C1 => n11689, C2 => 
                           n436, A => n14173, ZN => n14170);
   U12662 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_25_4_port, B1 => 
                           n458, B2 => REGISTERS_29_4_port, C1 => n469, C2 => 
                           REGISTERS_33_4_port, ZN => n14173);
   U12663 : OAI221_X1 port map( B1 => n11401, B2 => n480, C1 => n11529, C2 => 
                           n491, A => n14174, ZN => n14169);
   U12664 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_20_4_port, B1 => 
                           n513, B2 => REGISTERS_24_4_port, C1 => n524, C2 => 
                           REGISTERS_28_4_port, ZN => n14174);
   U12665 : OAI221_X1 port map( B1 => n11241, B2 => n535, C1 => n11369, C2 => 
                           n546, A => n14175, ZN => n14168);
   U12666 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_23_4_port, B1 => 
                           n568, B2 => REGISTERS_21_4_port, C1 => n579, C2 => 
                           REGISTERS_19_4_port, ZN => n14175);
   U12667 : NOR4_X1 port map( A1 => n14178, A2 => n14179, A3 => n14180, A4 => 
                           n14181, ZN => n14177);
   U12668 : OAI221_X1 port map( B1 => n11145, B2 => n315, C1 => n11081, C2 => 
                           n326, A => n14182, ZN => n14181);
   U12669 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_16_4_port, B1 => 
                           n119, B2 => REGISTERS_14_4_port, C1 => n13807, C2 =>
                           REGISTERS_12_4_port, ZN => n14182);
   U12670 : OAI221_X1 port map( B1 => n11113, B2 => n13863, C1 => n10857, C2 =>
                           n13809, A => n14183, ZN => n14180);
   U12671 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_4_port, B1 => 
                           n13865, B2 => REGISTERS_9_4_port, C1 => n13813, C2 
                           => REGISTERS_7_4_port, ZN => n14183);
   U12672 : OAI221_X1 port map( B1 => n10953, B2 => n13866, C1 => n10697, C2 =>
                           n13815, A => n14184, ZN => n14179);
   U12673 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_4_port, B1 => 
                           n13868, B2 => REGISTERS_36_4_port, C1 => n13819, C2 
                           => REGISTERS_3_4_port, ZN => n14184);
   U12674 : OAI221_X1 port map( B1 => n10793, B2 => n13869, C1 => n10665, C2 =>
                           n13821, A => n14185, ZN => n14178);
   U12675 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_4_port, B1 => 
                           n13871, B2 => REGISTERS_0_4_port, C1 => n13825, C2 
                           => REGISTERS_1_4_port, ZN => n14185);
   U12676 : NOR4_X1 port map( A1 => n14186, A2 => n14187, A3 => n14188, A4 => 
                           n14189, ZN => n14176);
   U12677 : OAI221_X1 port map( B1 => n11753, B2 => n370, C1 => n11017, C2 => 
                           n381, A => n14190, ZN => n14189);
   U12678 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_31_4_port, B1 => 
                           n403, B2 => REGISTERS_35_4_port, C1 => n414, C2 => 
                           REGISTERS_39_4_port, ZN => n14190);
   U12679 : OAI221_X1 port map( B1 => n11593, B2 => n425, C1 => n11721, C2 => 
                           n436, A => n14191, ZN => n14188);
   U12680 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_26_4_port, B1 => 
                           n458, B2 => REGISTERS_30_4_port, C1 => n469, C2 => 
                           REGISTERS_34_4_port, ZN => n14191);
   U12681 : OAI221_X1 port map( B1 => n11433, B2 => n480, C1 => n11561, C2 => 
                           n491, A => n14192, ZN => n14187);
   U12682 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_21_4_port, B1 => 
                           n513, B2 => REGISTERS_25_4_port, C1 => n524, C2 => 
                           REGISTERS_29_4_port, ZN => n14192);
   U12683 : OAI221_X1 port map( B1 => n11273, B2 => n535, C1 => n11401, C2 => 
                           n546, A => n14193, ZN => n14186);
   U12684 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_24_4_port, B1 => 
                           n568, B2 => REGISTERS_22_4_port, C1 => n579, C2 => 
                           REGISTERS_20_4_port, ZN => n14193);
   U12685 : AOI22_X1 port map( A1 => n13880, A2 => n4914, B1 => n13881, B2 => 
                           n4915, ZN => n14154);
   U12686 : NOR4_X1 port map( A1 => n14196, A2 => n14197, A3 => n14198, A4 => 
                           n14199, ZN => n14195);
   U12687 : OAI221_X1 port map( B1 => n11081, B2 => n315, C1 => n11017, C2 => 
                           n326, A => n14200, ZN => n14199);
   U12688 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_14_4_port, B1 => 
                           n13808, B2 => REGISTERS_38_4_port, C1 => n13889, C2 
                           => REGISTERS_39_4_port, ZN => n14200);
   U12689 : OAI221_X1 port map( B1 => n10921, B2 => n13810, C1 => n10857, C2 =>
                           n13890, A => n14201, ZN => n14198);
   U12690 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_4_port, B1 => 
                           n342, B2 => REGISTERS_9_4_port, C1 => n13812, C2 => 
                           REGISTERS_16_4_port, ZN => n14201);
   U12691 : OAI221_X1 port map( B1 => n10761, B2 => n303, C1 => n10697, C2 => 
                           n13893, A => n14202, ZN => n14197);
   U12692 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_4_port, B1 => 
                           n353, B2 => REGISTERS_4_4_port, C1 => n13818, C2 => 
                           REGISTERS_11_4_port, ZN => n14202);
   U12693 : OAI221_X1 port map( B1 => n11625, B2 => n304, C1 => n10569, C2 => 
                           n13896, A => n14203, ZN => n14196);
   U12694 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_4_port, B1 => 
                           n13826, B2 => REGISTERS_0_4_port, C1 => n13824, C2 
                           => REGISTERS_6_4_port, ZN => n14203);
   U12695 : NOR4_X1 port map( A1 => n14204, A2 => n14205, A3 => n14206, A4 => 
                           n14207, ZN => n14194);
   U12696 : OAI221_X1 port map( B1 => n11689, B2 => n370, C1 => n10953, C2 => 
                           n381, A => n14208, ZN => n14207);
   U12697 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_29_4_port, B1 => 
                           n403, B2 => REGISTERS_33_4_port, C1 => n414, C2 => 
                           REGISTERS_37_4_port, ZN => n14208);
   U12698 : OAI221_X1 port map( B1 => n11529, B2 => n425, C1 => n11657, C2 => 
                           n436, A => n14209, ZN => n14206);
   U12699 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_24_4_port, B1 => 
                           n458, B2 => REGISTERS_28_4_port, C1 => n469, C2 => 
                           REGISTERS_32_4_port, ZN => n14209);
   U12700 : OAI221_X1 port map( B1 => n11369, B2 => n480, C1 => n11497, C2 => 
                           n491, A => n14210, ZN => n14205);
   U12701 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_19_4_port, B1 => 
                           n513, B2 => REGISTERS_23_4_port, C1 => n524, C2 => 
                           REGISTERS_27_4_port, ZN => n14210);
   U12702 : OAI221_X1 port map( B1 => n11209, B2 => n535, C1 => n11337, C2 => 
                           n546, A => n14211, ZN => n14204);
   U12703 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_22_4_port, B1 => 
                           n568, B2 => REGISTERS_20_4_port, C1 => n579, C2 => 
                           REGISTERS_18_4_port, ZN => n14211);
   U12704 : NOR4_X1 port map( A1 => n14214, A2 => n14215, A3 => n14216, A4 => 
                           n14217, ZN => n14213);
   U12705 : OAI221_X1 port map( B1 => n11049, B2 => n315, C1 => n10985, C2 => 
                           n326, A => n14218, ZN => n14217);
   U12706 : AOI222_X1 port map( A1 => n337, A2 => REGISTERS_13_4_port, B1 => 
                           n13808, B2 => REGISTERS_37_4_port, C1 => n13889, C2 
                           => REGISTERS_38_4_port, ZN => n14218);
   U12707 : OAI221_X1 port map( B1 => n10889, B2 => n13810, C1 => n10825, C2 =>
                           n13890, A => n14219, ZN => n14216);
   U12708 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_4_port, B1 => 
                           n342, B2 => REGISTERS_8_4_port, C1 => n13812, C2 => 
                           REGISTERS_15_4_port, ZN => n14219);
   U12709 : OAI221_X1 port map( B1 => n10729, B2 => n303, C1 => n10665, C2 => 
                           n13893, A => n14220, ZN => n14215);
   U12710 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_4_port, B1 => 
                           n353, B2 => REGISTERS_3_4_port, C1 => n13818, C2 => 
                           REGISTERS_10_4_port, ZN => n14220);
   U12711 : OAI221_X1 port map( B1 => n11593, B2 => n304, C1 => n10529, C2 => 
                           n13896, A => n14221, ZN => n14214);
   U12712 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_4_port, B1 => 
                           n13917, B2 => REGISTERS_39_4_port, C1 => n13824, C2 
                           => REGISTERS_5_4_port, ZN => n14221);
   U12713 : NOR4_X1 port map( A1 => n14222, A2 => n14223, A3 => n14224, A4 => 
                           n14225, ZN => n14212);
   U12714 : OAI221_X1 port map( B1 => n11657, B2 => n370, C1 => n10921, C2 => 
                           n381, A => n14226, ZN => n14225);
   U12715 : AOI222_X1 port map( A1 => n392, A2 => REGISTERS_28_4_port, B1 => 
                           n403, B2 => REGISTERS_32_4_port, C1 => n414, C2 => 
                           REGISTERS_36_4_port, ZN => n14226);
   U12716 : OAI221_X1 port map( B1 => n11497, B2 => n425, C1 => n11625, C2 => 
                           n436, A => n14227, ZN => n14224);
   U12717 : AOI222_X1 port map( A1 => n447, A2 => REGISTERS_23_4_port, B1 => 
                           n458, B2 => REGISTERS_27_4_port, C1 => n469, C2 => 
                           REGISTERS_31_4_port, ZN => n14227);
   U12718 : OAI221_X1 port map( B1 => n11337, B2 => n480, C1 => n11465, C2 => 
                           n491, A => n14228, ZN => n14223);
   U12719 : AOI222_X1 port map( A1 => n502, A2 => REGISTERS_18_4_port, B1 => 
                           n513, B2 => REGISTERS_22_4_port, C1 => n524, C2 => 
                           REGISTERS_26_4_port, ZN => n14228);
   U12720 : OAI221_X1 port map( B1 => n11177, B2 => n535, C1 => n11305, C2 => 
                           n546, A => n14229, ZN => n14222);
   U12721 : AOI222_X1 port map( A1 => n557, A2 => REGISTERS_21_4_port, B1 => 
                           n568, B2 => REGISTERS_19_4_port, C1 => n579, C2 => 
                           REGISTERS_17_4_port, ZN => n14229);
   U12722 : NAND3_X1 port map( A1 => n14230, A2 => n14231, A3 => n14232, ZN => 
                           n11899);
   U12723 : AOI221_X1 port map( B1 => n13792, B2 => n4919, C1 => n13793, C2 => 
                           MEM_IN(5), A => n14233, ZN => n14232);
   U12724 : OAI22_X1 port map( A1 => n10526, A2 => n251, B1 => n4921, B2 => 
                           n121, ZN => n14233);
   U12725 : NOR2_X1 port map( A1 => n5571, A2 => n13796, ZN => n5569);
   U12726 : INV_X1 port map( A => MEM_IN(5), ZN => n5571);
   U12727 : AOI22_X1 port map( A1 => n197, A2 => n4922, B1 => n150, B2 => n4923
                           , ZN => n14231);
   U12728 : NOR4_X1 port map( A1 => n14236, A2 => n14237, A3 => n14238, A4 => 
                           n14239, ZN => n14235);
   U12729 : OAI221_X1 port map( B1 => n11112, B2 => n314, C1 => n11048, C2 => 
                           n325, A => n14240, ZN => n14239);
   U12730 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_15_5_port, B1 => 
                           n13807, B2 => REGISTERS_11_5_port, C1 => n13808, C2 
                           => REGISTERS_39_5_port, ZN => n14240);
   U12731 : OAI221_X1 port map( B1 => n10824, B2 => n13809, C1 => n10952, C2 =>
                           n13810, A => n14241, ZN => n14238);
   U12732 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_5_port, B1 => 
                           n13813, B2 => REGISTERS_6_5_port, C1 => n347, C2 => 
                           REGISTERS_10_5_port, ZN => n14241);
   U12733 : OAI221_X1 port map( B1 => n10664, B2 => n13815, C1 => n10792, C2 =>
                           n303, A => n14242, ZN => n14237);
   U12734 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_5_port, B1 => 
                           n13819, B2 => REGISTERS_2_5_port, C1 => n358, C2 => 
                           REGISTERS_5_5_port, ZN => n14242);
   U12735 : OAI221_X1 port map( B1 => n10632, B2 => n13821, C1 => n11656, C2 =>
                           n304, A => n14243, ZN => n14236);
   U12736 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_5_port, B1 => 
                           n13825, B2 => REGISTERS_0_5_port, C1 => n13826, C2 
                           => REGISTERS_1_5_port, ZN => n14243);
   U12737 : NOR4_X1 port map( A1 => n14244, A2 => n14245, A3 => n14246, A4 => 
                           n14247, ZN => n14234);
   U12738 : OAI221_X1 port map( B1 => n11720, B2 => n369, C1 => n10984, C2 => 
                           n381, A => n14248, ZN => n14247);
   U12739 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_30_5_port, B1 => 
                           n402, B2 => REGISTERS_34_5_port, C1 => n413, C2 => 
                           REGISTERS_38_5_port, ZN => n14248);
   U12740 : OAI221_X1 port map( B1 => n11560, B2 => n424, C1 => n11688, C2 => 
                           n435, A => n14249, ZN => n14246);
   U12741 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_25_5_port, B1 => 
                           n457, B2 => REGISTERS_29_5_port, C1 => n468, C2 => 
                           REGISTERS_33_5_port, ZN => n14249);
   U12742 : OAI221_X1 port map( B1 => n11400, B2 => n479, C1 => n11528, C2 => 
                           n490, A => n14250, ZN => n14245);
   U12743 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_20_5_port, B1 => 
                           n512, B2 => REGISTERS_24_5_port, C1 => n523, C2 => 
                           REGISTERS_28_5_port, ZN => n14250);
   U12744 : OAI221_X1 port map( B1 => n11240, B2 => n534, C1 => n11368, C2 => 
                           n545, A => n14251, ZN => n14244);
   U12745 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_23_5_port, B1 => 
                           n567, B2 => REGISTERS_21_5_port, C1 => n578, C2 => 
                           REGISTERS_19_5_port, ZN => n14251);
   U12746 : NOR4_X1 port map( A1 => n14254, A2 => n14255, A3 => n14256, A4 => 
                           n14257, ZN => n14253);
   U12747 : OAI221_X1 port map( B1 => n11144, B2 => n314, C1 => n11080, C2 => 
                           n325, A => n14258, ZN => n14257);
   U12748 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_16_5_port, B1 => 
                           n119, B2 => REGISTERS_14_5_port, C1 => n13807, C2 =>
                           REGISTERS_12_5_port, ZN => n14258);
   U12749 : OAI221_X1 port map( B1 => n11112, B2 => n13863, C1 => n10856, C2 =>
                           n13809, A => n14259, ZN => n14256);
   U12750 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_5_port, B1 => 
                           n13865, B2 => REGISTERS_9_5_port, C1 => n13813, C2 
                           => REGISTERS_7_5_port, ZN => n14259);
   U12751 : OAI221_X1 port map( B1 => n10952, B2 => n13866, C1 => n10696, C2 =>
                           n13815, A => n14260, ZN => n14255);
   U12752 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_5_port, B1 => 
                           n13868, B2 => REGISTERS_36_5_port, C1 => n13819, C2 
                           => REGISTERS_3_5_port, ZN => n14260);
   U12753 : OAI221_X1 port map( B1 => n10792, B2 => n13869, C1 => n10664, C2 =>
                           n13821, A => n14261, ZN => n14254);
   U12754 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_5_port, B1 => 
                           n13871, B2 => REGISTERS_0_5_port, C1 => n13825, C2 
                           => REGISTERS_1_5_port, ZN => n14261);
   U12755 : NOR4_X1 port map( A1 => n14262, A2 => n14263, A3 => n14264, A4 => 
                           n14265, ZN => n14252);
   U12756 : OAI221_X1 port map( B1 => n11752, B2 => n369, C1 => n11016, C2 => 
                           n380, A => n14266, ZN => n14265);
   U12757 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_31_5_port, B1 => 
                           n402, B2 => REGISTERS_35_5_port, C1 => n413, C2 => 
                           REGISTERS_39_5_port, ZN => n14266);
   U12758 : OAI221_X1 port map( B1 => n11592, B2 => n424, C1 => n11720, C2 => 
                           n435, A => n14267, ZN => n14264);
   U12759 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_26_5_port, B1 => 
                           n457, B2 => REGISTERS_30_5_port, C1 => n468, C2 => 
                           REGISTERS_34_5_port, ZN => n14267);
   U12760 : OAI221_X1 port map( B1 => n11432, B2 => n479, C1 => n11560, C2 => 
                           n490, A => n14268, ZN => n14263);
   U12761 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_21_5_port, B1 => 
                           n512, B2 => REGISTERS_25_5_port, C1 => n523, C2 => 
                           REGISTERS_29_5_port, ZN => n14268);
   U12762 : OAI221_X1 port map( B1 => n11272, B2 => n534, C1 => n11400, C2 => 
                           n545, A => n14269, ZN => n14262);
   U12763 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_24_5_port, B1 => 
                           n567, B2 => REGISTERS_22_5_port, C1 => n578, C2 => 
                           REGISTERS_20_5_port, ZN => n14269);
   U12764 : AOI22_X1 port map( A1 => n13880, A2 => n4924, B1 => n13881, B2 => 
                           n4925, ZN => n14230);
   U12765 : NOR4_X1 port map( A1 => n14272, A2 => n14273, A3 => n14274, A4 => 
                           n14275, ZN => n14271);
   U12766 : OAI221_X1 port map( B1 => n11080, B2 => n314, C1 => n11016, C2 => 
                           n325, A => n14276, ZN => n14275);
   U12767 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_14_5_port, B1 => 
                           n13808, B2 => REGISTERS_38_5_port, C1 => n13889, C2 
                           => REGISTERS_39_5_port, ZN => n14276);
   U12768 : OAI221_X1 port map( B1 => n10920, B2 => n13810, C1 => n10856, C2 =>
                           n13890, A => n14277, ZN => n14274);
   U12769 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_5_port, B1 => 
                           n341, B2 => REGISTERS_9_5_port, C1 => n13812, C2 => 
                           REGISTERS_16_5_port, ZN => n14277);
   U12770 : OAI221_X1 port map( B1 => n10760, B2 => n303, C1 => n10696, C2 => 
                           n13893, A => n14278, ZN => n14273);
   U12771 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_5_port, B1 => 
                           n352, B2 => REGISTERS_4_5_port, C1 => n13818, C2 => 
                           REGISTERS_11_5_port, ZN => n14278);
   U12772 : OAI221_X1 port map( B1 => n11624, B2 => n304, C1 => n10568, C2 => 
                           n13896, A => n14279, ZN => n14272);
   U12773 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_5_port, B1 => 
                           n13826, B2 => REGISTERS_0_5_port, C1 => n13824, C2 
                           => REGISTERS_6_5_port, ZN => n14279);
   U12774 : NOR4_X1 port map( A1 => n14280, A2 => n14281, A3 => n14282, A4 => 
                           n14283, ZN => n14270);
   U12775 : OAI221_X1 port map( B1 => n11688, B2 => n369, C1 => n10952, C2 => 
                           n380, A => n14284, ZN => n14283);
   U12776 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_29_5_port, B1 => 
                           n402, B2 => REGISTERS_33_5_port, C1 => n413, C2 => 
                           REGISTERS_37_5_port, ZN => n14284);
   U12777 : OAI221_X1 port map( B1 => n11528, B2 => n424, C1 => n11656, C2 => 
                           n435, A => n14285, ZN => n14282);
   U12778 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_24_5_port, B1 => 
                           n457, B2 => REGISTERS_28_5_port, C1 => n468, C2 => 
                           REGISTERS_32_5_port, ZN => n14285);
   U12779 : OAI221_X1 port map( B1 => n11368, B2 => n479, C1 => n11496, C2 => 
                           n490, A => n14286, ZN => n14281);
   U12780 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_19_5_port, B1 => 
                           n512, B2 => REGISTERS_23_5_port, C1 => n523, C2 => 
                           REGISTERS_27_5_port, ZN => n14286);
   U12781 : OAI221_X1 port map( B1 => n11208, B2 => n534, C1 => n11336, C2 => 
                           n545, A => n14287, ZN => n14280);
   U12782 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_22_5_port, B1 => 
                           n567, B2 => REGISTERS_20_5_port, C1 => n578, C2 => 
                           REGISTERS_18_5_port, ZN => n14287);
   U12783 : NOR4_X1 port map( A1 => n14290, A2 => n14291, A3 => n14292, A4 => 
                           n14293, ZN => n14289);
   U12784 : OAI221_X1 port map( B1 => n11048, B2 => n314, C1 => n10984, C2 => 
                           n325, A => n14294, ZN => n14293);
   U12785 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_13_5_port, B1 => 
                           n13808, B2 => REGISTERS_37_5_port, C1 => n13889, C2 
                           => REGISTERS_38_5_port, ZN => n14294);
   U12786 : OAI221_X1 port map( B1 => n10888, B2 => n13810, C1 => n10824, C2 =>
                           n13890, A => n14295, ZN => n14292);
   U12787 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_5_port, B1 => 
                           n342, B2 => REGISTERS_8_5_port, C1 => n13812, C2 => 
                           REGISTERS_15_5_port, ZN => n14295);
   U12788 : OAI221_X1 port map( B1 => n10728, B2 => n303, C1 => n10664, C2 => 
                           n13893, A => n14296, ZN => n14291);
   U12789 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_5_port, B1 => 
                           n353, B2 => REGISTERS_3_5_port, C1 => n13818, C2 => 
                           REGISTERS_10_5_port, ZN => n14296);
   U12790 : OAI221_X1 port map( B1 => n11592, B2 => n304, C1 => n10526, C2 => 
                           n13896, A => n14297, ZN => n14290);
   U12791 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_5_port, B1 => 
                           n13917, B2 => REGISTERS_39_5_port, C1 => n13824, C2 
                           => REGISTERS_5_5_port, ZN => n14297);
   U12792 : NOR4_X1 port map( A1 => n14298, A2 => n14299, A3 => n14300, A4 => 
                           n14301, ZN => n14288);
   U12793 : OAI221_X1 port map( B1 => n11656, B2 => n369, C1 => n10920, C2 => 
                           n380, A => n14302, ZN => n14301);
   U12794 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_28_5_port, B1 => 
                           n402, B2 => REGISTERS_32_5_port, C1 => n413, C2 => 
                           REGISTERS_36_5_port, ZN => n14302);
   U12795 : OAI221_X1 port map( B1 => n11496, B2 => n424, C1 => n11624, C2 => 
                           n435, A => n14303, ZN => n14300);
   U12796 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_23_5_port, B1 => 
                           n457, B2 => REGISTERS_27_5_port, C1 => n468, C2 => 
                           REGISTERS_31_5_port, ZN => n14303);
   U12797 : OAI221_X1 port map( B1 => n11336, B2 => n479, C1 => n11464, C2 => 
                           n490, A => n14304, ZN => n14299);
   U12798 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_18_5_port, B1 => 
                           n512, B2 => REGISTERS_22_5_port, C1 => n523, C2 => 
                           REGISTERS_26_5_port, ZN => n14304);
   U12799 : OAI221_X1 port map( B1 => n11176, B2 => n534, C1 => n11304, C2 => 
                           n545, A => n14305, ZN => n14298);
   U12800 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_21_5_port, B1 => 
                           n567, B2 => REGISTERS_19_5_port, C1 => n578, C2 => 
                           REGISTERS_17_5_port, ZN => n14305);
   U12801 : NAND3_X1 port map( A1 => n14306, A2 => n14307, A3 => n14308, ZN => 
                           n11898);
   U12802 : AOI221_X1 port map( B1 => n13792, B2 => n4929, C1 => n13793, C2 => 
                           MEM_IN(6), A => n14309, ZN => n14308);
   U12803 : OAI22_X1 port map( A1 => n10523, A2 => n251, B1 => n4931, B2 => 
                           n121, ZN => n14309);
   U12804 : NOR2_X1 port map( A1 => n5578, A2 => n13796, ZN => n5576);
   U12805 : INV_X1 port map( A => MEM_IN(6), ZN => n5578);
   U12806 : AOI22_X1 port map( A1 => n197, A2 => n4932, B1 => n150, B2 => n4933
                           , ZN => n14307);
   U12807 : NOR4_X1 port map( A1 => n14312, A2 => n14313, A3 => n14314, A4 => 
                           n14315, ZN => n14311);
   U12808 : OAI221_X1 port map( B1 => n11111, B2 => n314, C1 => n11047, C2 => 
                           n325, A => n14316, ZN => n14315);
   U12809 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_15_6_port, B1 => 
                           n13807, B2 => REGISTERS_11_6_port, C1 => n13808, C2 
                           => REGISTERS_39_6_port, ZN => n14316);
   U12810 : OAI221_X1 port map( B1 => n10823, B2 => n13809, C1 => n10951, C2 =>
                           n13810, A => n14317, ZN => n14314);
   U12811 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_6_port, B1 => 
                           n13813, B2 => REGISTERS_6_6_port, C1 => n347, C2 => 
                           REGISTERS_10_6_port, ZN => n14317);
   U12812 : OAI221_X1 port map( B1 => n10663, B2 => n13815, C1 => n10791, C2 =>
                           n303, A => n14318, ZN => n14313);
   U12813 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_6_port, B1 => 
                           n13819, B2 => REGISTERS_2_6_port, C1 => n358, C2 => 
                           REGISTERS_5_6_port, ZN => n14318);
   U12814 : OAI221_X1 port map( B1 => n10631, B2 => n13821, C1 => n11655, C2 =>
                           n304, A => n14319, ZN => n14312);
   U12815 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_6_port, B1 => 
                           n13825, B2 => REGISTERS_0_6_port, C1 => n13826, C2 
                           => REGISTERS_1_6_port, ZN => n14319);
   U12816 : NOR4_X1 port map( A1 => n14320, A2 => n14321, A3 => n14322, A4 => 
                           n14323, ZN => n14310);
   U12817 : OAI221_X1 port map( B1 => n11719, B2 => n369, C1 => n10983, C2 => 
                           n380, A => n14324, ZN => n14323);
   U12818 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_30_6_port, B1 => 
                           n402, B2 => REGISTERS_34_6_port, C1 => n413, C2 => 
                           REGISTERS_38_6_port, ZN => n14324);
   U12819 : OAI221_X1 port map( B1 => n11559, B2 => n424, C1 => n11687, C2 => 
                           n435, A => n14325, ZN => n14322);
   U12820 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_25_6_port, B1 => 
                           n457, B2 => REGISTERS_29_6_port, C1 => n468, C2 => 
                           REGISTERS_33_6_port, ZN => n14325);
   U12821 : OAI221_X1 port map( B1 => n11399, B2 => n479, C1 => n11527, C2 => 
                           n490, A => n14326, ZN => n14321);
   U12822 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_20_6_port, B1 => 
                           n512, B2 => REGISTERS_24_6_port, C1 => n523, C2 => 
                           REGISTERS_28_6_port, ZN => n14326);
   U12823 : OAI221_X1 port map( B1 => n11239, B2 => n534, C1 => n11367, C2 => 
                           n545, A => n14327, ZN => n14320);
   U12824 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_23_6_port, B1 => 
                           n567, B2 => REGISTERS_21_6_port, C1 => n578, C2 => 
                           REGISTERS_19_6_port, ZN => n14327);
   U12825 : NOR4_X1 port map( A1 => n14330, A2 => n14331, A3 => n14332, A4 => 
                           n14333, ZN => n14329);
   U12826 : OAI221_X1 port map( B1 => n11143, B2 => n314, C1 => n11079, C2 => 
                           n325, A => n14334, ZN => n14333);
   U12827 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_16_6_port, B1 => 
                           n119, B2 => REGISTERS_14_6_port, C1 => n13807, C2 =>
                           REGISTERS_12_6_port, ZN => n14334);
   U12828 : OAI221_X1 port map( B1 => n11111, B2 => n13863, C1 => n10855, C2 =>
                           n13809, A => n14335, ZN => n14332);
   U12829 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_6_port, B1 => 
                           n13865, B2 => REGISTERS_9_6_port, C1 => n13813, C2 
                           => REGISTERS_7_6_port, ZN => n14335);
   U12830 : OAI221_X1 port map( B1 => n10951, B2 => n13866, C1 => n10695, C2 =>
                           n13815, A => n14336, ZN => n14331);
   U12831 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_6_port, B1 => 
                           n13868, B2 => REGISTERS_36_6_port, C1 => n13819, C2 
                           => REGISTERS_3_6_port, ZN => n14336);
   U12832 : OAI221_X1 port map( B1 => n10791, B2 => n13869, C1 => n10663, C2 =>
                           n13821, A => n14337, ZN => n14330);
   U12833 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_6_port, B1 => 
                           n13871, B2 => REGISTERS_0_6_port, C1 => n13825, C2 
                           => REGISTERS_1_6_port, ZN => n14337);
   U12834 : NOR4_X1 port map( A1 => n14338, A2 => n14339, A3 => n14340, A4 => 
                           n14341, ZN => n14328);
   U12835 : OAI221_X1 port map( B1 => n11751, B2 => n369, C1 => n11015, C2 => 
                           n380, A => n14342, ZN => n14341);
   U12836 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_31_6_port, B1 => 
                           n402, B2 => REGISTERS_35_6_port, C1 => n413, C2 => 
                           REGISTERS_39_6_port, ZN => n14342);
   U12837 : OAI221_X1 port map( B1 => n11591, B2 => n424, C1 => n11719, C2 => 
                           n435, A => n14343, ZN => n14340);
   U12838 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_26_6_port, B1 => 
                           n457, B2 => REGISTERS_30_6_port, C1 => n468, C2 => 
                           REGISTERS_34_6_port, ZN => n14343);
   U12839 : OAI221_X1 port map( B1 => n11431, B2 => n479, C1 => n11559, C2 => 
                           n490, A => n14344, ZN => n14339);
   U12840 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_21_6_port, B1 => 
                           n512, B2 => REGISTERS_25_6_port, C1 => n523, C2 => 
                           REGISTERS_29_6_port, ZN => n14344);
   U12841 : OAI221_X1 port map( B1 => n11271, B2 => n534, C1 => n11399, C2 => 
                           n545, A => n14345, ZN => n14338);
   U12842 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_24_6_port, B1 => 
                           n567, B2 => REGISTERS_22_6_port, C1 => n578, C2 => 
                           REGISTERS_20_6_port, ZN => n14345);
   U12843 : AOI22_X1 port map( A1 => n13880, A2 => n4934, B1 => n13881, B2 => 
                           n4935, ZN => n14306);
   U12844 : NOR4_X1 port map( A1 => n14348, A2 => n14349, A3 => n14350, A4 => 
                           n14351, ZN => n14347);
   U12845 : OAI221_X1 port map( B1 => n11079, B2 => n314, C1 => n11015, C2 => 
                           n325, A => n14352, ZN => n14351);
   U12846 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_14_6_port, B1 => 
                           n13808, B2 => REGISTERS_38_6_port, C1 => n13889, C2 
                           => REGISTERS_39_6_port, ZN => n14352);
   U12847 : OAI221_X1 port map( B1 => n10919, B2 => n13810, C1 => n10855, C2 =>
                           n13890, A => n14353, ZN => n14350);
   U12848 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_6_port, B1 => 
                           n342, B2 => REGISTERS_9_6_port, C1 => n13812, C2 => 
                           REGISTERS_16_6_port, ZN => n14353);
   U12849 : OAI221_X1 port map( B1 => n10759, B2 => n303, C1 => n10695, C2 => 
                           n13893, A => n14354, ZN => n14349);
   U12850 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_6_port, B1 => 
                           n353, B2 => REGISTERS_4_6_port, C1 => n13818, C2 => 
                           REGISTERS_11_6_port, ZN => n14354);
   U12851 : OAI221_X1 port map( B1 => n11623, B2 => n304, C1 => n10567, C2 => 
                           n13896, A => n14355, ZN => n14348);
   U12852 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_6_port, B1 => 
                           n13826, B2 => REGISTERS_0_6_port, C1 => n13824, C2 
                           => REGISTERS_6_6_port, ZN => n14355);
   U12853 : NOR4_X1 port map( A1 => n14356, A2 => n14357, A3 => n14358, A4 => 
                           n14359, ZN => n14346);
   U12854 : OAI221_X1 port map( B1 => n11687, B2 => n369, C1 => n10951, C2 => 
                           n380, A => n14360, ZN => n14359);
   U12855 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_29_6_port, B1 => 
                           n402, B2 => REGISTERS_33_6_port, C1 => n413, C2 => 
                           REGISTERS_37_6_port, ZN => n14360);
   U12856 : OAI221_X1 port map( B1 => n11527, B2 => n424, C1 => n11655, C2 => 
                           n435, A => n14361, ZN => n14358);
   U12857 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_24_6_port, B1 => 
                           n457, B2 => REGISTERS_28_6_port, C1 => n468, C2 => 
                           REGISTERS_32_6_port, ZN => n14361);
   U12858 : OAI221_X1 port map( B1 => n11367, B2 => n479, C1 => n11495, C2 => 
                           n490, A => n14362, ZN => n14357);
   U12859 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_19_6_port, B1 => 
                           n512, B2 => REGISTERS_23_6_port, C1 => n523, C2 => 
                           REGISTERS_27_6_port, ZN => n14362);
   U12860 : OAI221_X1 port map( B1 => n11207, B2 => n534, C1 => n11335, C2 => 
                           n545, A => n14363, ZN => n14356);
   U12861 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_22_6_port, B1 => 
                           n567, B2 => REGISTERS_20_6_port, C1 => n578, C2 => 
                           REGISTERS_18_6_port, ZN => n14363);
   U12862 : NOR4_X1 port map( A1 => n14366, A2 => n14367, A3 => n14368, A4 => 
                           n14369, ZN => n14365);
   U12863 : OAI221_X1 port map( B1 => n11047, B2 => n314, C1 => n10983, C2 => 
                           n325, A => n14370, ZN => n14369);
   U12864 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_13_6_port, B1 => 
                           n13808, B2 => REGISTERS_37_6_port, C1 => n13889, C2 
                           => REGISTERS_38_6_port, ZN => n14370);
   U12865 : OAI221_X1 port map( B1 => n10887, B2 => n13810, C1 => n10823, C2 =>
                           n13890, A => n14371, ZN => n14368);
   U12866 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_6_port, B1 => 
                           n342, B2 => REGISTERS_8_6_port, C1 => n13812, C2 => 
                           REGISTERS_15_6_port, ZN => n14371);
   U12867 : OAI221_X1 port map( B1 => n10727, B2 => n303, C1 => n10663, C2 => 
                           n13893, A => n14372, ZN => n14367);
   U12868 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_6_port, B1 => 
                           n353, B2 => REGISTERS_3_6_port, C1 => n13818, C2 => 
                           REGISTERS_10_6_port, ZN => n14372);
   U12869 : OAI221_X1 port map( B1 => n11591, B2 => n304, C1 => n10523, C2 => 
                           n13896, A => n14373, ZN => n14366);
   U12870 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_6_port, B1 => 
                           n13917, B2 => REGISTERS_39_6_port, C1 => n13824, C2 
                           => REGISTERS_5_6_port, ZN => n14373);
   U12871 : NOR4_X1 port map( A1 => n14374, A2 => n14375, A3 => n14376, A4 => 
                           n14377, ZN => n14364);
   U12872 : OAI221_X1 port map( B1 => n11655, B2 => n369, C1 => n10919, C2 => 
                           n380, A => n14378, ZN => n14377);
   U12873 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_28_6_port, B1 => 
                           n402, B2 => REGISTERS_32_6_port, C1 => n413, C2 => 
                           REGISTERS_36_6_port, ZN => n14378);
   U12874 : OAI221_X1 port map( B1 => n11495, B2 => n424, C1 => n11623, C2 => 
                           n435, A => n14379, ZN => n14376);
   U12875 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_23_6_port, B1 => 
                           n457, B2 => REGISTERS_27_6_port, C1 => n468, C2 => 
                           REGISTERS_31_6_port, ZN => n14379);
   U12876 : OAI221_X1 port map( B1 => n11335, B2 => n479, C1 => n11463, C2 => 
                           n490, A => n14380, ZN => n14375);
   U12877 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_18_6_port, B1 => 
                           n512, B2 => REGISTERS_22_6_port, C1 => n523, C2 => 
                           REGISTERS_26_6_port, ZN => n14380);
   U12878 : OAI221_X1 port map( B1 => n11175, B2 => n534, C1 => n11303, C2 => 
                           n545, A => n14381, ZN => n14374);
   U12879 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_21_6_port, B1 => 
                           n567, B2 => REGISTERS_19_6_port, C1 => n578, C2 => 
                           REGISTERS_17_6_port, ZN => n14381);
   U12880 : NAND3_X1 port map( A1 => n14382, A2 => n14383, A3 => n14384, ZN => 
                           n11897);
   U12881 : AOI221_X1 port map( B1 => n13792, B2 => n4939, C1 => n13793, C2 => 
                           MEM_IN(7), A => n14385, ZN => n14384);
   U12882 : OAI22_X1 port map( A1 => n10520, A2 => n251, B1 => n4941, B2 => 
                           n121, ZN => n14385);
   U12883 : NOR2_X1 port map( A1 => n5585, A2 => n13796, ZN => n5583);
   U12884 : INV_X1 port map( A => MEM_IN(7), ZN => n5585);
   U12885 : AOI22_X1 port map( A1 => n197, A2 => n4942, B1 => n150, B2 => n4943
                           , ZN => n14383);
   U12886 : NOR4_X1 port map( A1 => n14388, A2 => n14389, A3 => n14390, A4 => 
                           n14391, ZN => n14387);
   U12887 : OAI221_X1 port map( B1 => n11110, B2 => n314, C1 => n11046, C2 => 
                           n325, A => n14392, ZN => n14391);
   U12888 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_15_7_port, B1 => 
                           n13807, B2 => REGISTERS_11_7_port, C1 => n13808, C2 
                           => REGISTERS_39_7_port, ZN => n14392);
   U12889 : OAI221_X1 port map( B1 => n10822, B2 => n13809, C1 => n10950, C2 =>
                           n13810, A => n14393, ZN => n14390);
   U12890 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_7_port, B1 => 
                           n13813, B2 => REGISTERS_6_7_port, C1 => n347, C2 => 
                           REGISTERS_10_7_port, ZN => n14393);
   U12891 : OAI221_X1 port map( B1 => n10662, B2 => n13815, C1 => n10790, C2 =>
                           n303, A => n14394, ZN => n14389);
   U12892 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_7_port, B1 => 
                           n13819, B2 => REGISTERS_2_7_port, C1 => n358, C2 => 
                           REGISTERS_5_7_port, ZN => n14394);
   U12893 : OAI221_X1 port map( B1 => n10630, B2 => n13821, C1 => n11654, C2 =>
                           n304, A => n14395, ZN => n14388);
   U12894 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_7_port, B1 => 
                           n13825, B2 => REGISTERS_0_7_port, C1 => n13826, C2 
                           => REGISTERS_1_7_port, ZN => n14395);
   U12895 : NOR4_X1 port map( A1 => n14396, A2 => n14397, A3 => n14398, A4 => 
                           n14399, ZN => n14386);
   U12896 : OAI221_X1 port map( B1 => n11718, B2 => n369, C1 => n10982, C2 => 
                           n380, A => n14400, ZN => n14399);
   U12897 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_30_7_port, B1 => 
                           n402, B2 => REGISTERS_34_7_port, C1 => n413, C2 => 
                           REGISTERS_38_7_port, ZN => n14400);
   U12898 : OAI221_X1 port map( B1 => n11558, B2 => n424, C1 => n11686, C2 => 
                           n435, A => n14401, ZN => n14398);
   U12899 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_25_7_port, B1 => 
                           n457, B2 => REGISTERS_29_7_port, C1 => n468, C2 => 
                           REGISTERS_33_7_port, ZN => n14401);
   U12900 : OAI221_X1 port map( B1 => n11398, B2 => n479, C1 => n11526, C2 => 
                           n490, A => n14402, ZN => n14397);
   U12901 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_20_7_port, B1 => 
                           n512, B2 => REGISTERS_24_7_port, C1 => n523, C2 => 
                           REGISTERS_28_7_port, ZN => n14402);
   U12902 : OAI221_X1 port map( B1 => n11238, B2 => n534, C1 => n11366, C2 => 
                           n545, A => n14403, ZN => n14396);
   U12903 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_23_7_port, B1 => 
                           n567, B2 => REGISTERS_21_7_port, C1 => n578, C2 => 
                           REGISTERS_19_7_port, ZN => n14403);
   U12904 : NOR4_X1 port map( A1 => n14406, A2 => n14407, A3 => n14408, A4 => 
                           n14409, ZN => n14405);
   U12905 : OAI221_X1 port map( B1 => n11142, B2 => n314, C1 => n11078, C2 => 
                           n325, A => n14410, ZN => n14409);
   U12906 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_16_7_port, B1 => 
                           n119, B2 => REGISTERS_14_7_port, C1 => n13807, C2 =>
                           REGISTERS_12_7_port, ZN => n14410);
   U12907 : OAI221_X1 port map( B1 => n11110, B2 => n13863, C1 => n10854, C2 =>
                           n13809, A => n14411, ZN => n14408);
   U12908 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_7_port, B1 => 
                           n13865, B2 => REGISTERS_9_7_port, C1 => n13813, C2 
                           => REGISTERS_7_7_port, ZN => n14411);
   U12909 : OAI221_X1 port map( B1 => n10950, B2 => n13866, C1 => n10694, C2 =>
                           n13815, A => n14412, ZN => n14407);
   U12910 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_7_port, B1 => 
                           n13868, B2 => REGISTERS_36_7_port, C1 => n13819, C2 
                           => REGISTERS_3_7_port, ZN => n14412);
   U12911 : OAI221_X1 port map( B1 => n10790, B2 => n13869, C1 => n10662, C2 =>
                           n13821, A => n14413, ZN => n14406);
   U12912 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_7_port, B1 => 
                           n13871, B2 => REGISTERS_0_7_port, C1 => n13825, C2 
                           => REGISTERS_1_7_port, ZN => n14413);
   U12913 : NOR4_X1 port map( A1 => n14414, A2 => n14415, A3 => n14416, A4 => 
                           n14417, ZN => n14404);
   U12914 : OAI221_X1 port map( B1 => n11750, B2 => n369, C1 => n11014, C2 => 
                           n380, A => n14418, ZN => n14417);
   U12915 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_31_7_port, B1 => 
                           n402, B2 => REGISTERS_35_7_port, C1 => n413, C2 => 
                           REGISTERS_39_7_port, ZN => n14418);
   U12916 : OAI221_X1 port map( B1 => n11590, B2 => n424, C1 => n11718, C2 => 
                           n435, A => n14419, ZN => n14416);
   U12917 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_26_7_port, B1 => 
                           n457, B2 => REGISTERS_30_7_port, C1 => n468, C2 => 
                           REGISTERS_34_7_port, ZN => n14419);
   U12918 : OAI221_X1 port map( B1 => n11430, B2 => n479, C1 => n11558, C2 => 
                           n490, A => n14420, ZN => n14415);
   U12919 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_21_7_port, B1 => 
                           n512, B2 => REGISTERS_25_7_port, C1 => n523, C2 => 
                           REGISTERS_29_7_port, ZN => n14420);
   U12920 : OAI221_X1 port map( B1 => n11270, B2 => n534, C1 => n11398, C2 => 
                           n545, A => n14421, ZN => n14414);
   U12921 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_24_7_port, B1 => 
                           n567, B2 => REGISTERS_22_7_port, C1 => n578, C2 => 
                           REGISTERS_20_7_port, ZN => n14421);
   U12922 : AOI22_X1 port map( A1 => n13880, A2 => n4944, B1 => n13881, B2 => 
                           n4945, ZN => n14382);
   U12923 : NOR4_X1 port map( A1 => n14424, A2 => n14425, A3 => n14426, A4 => 
                           n14427, ZN => n14423);
   U12924 : OAI221_X1 port map( B1 => n11078, B2 => n314, C1 => n11014, C2 => 
                           n325, A => n14428, ZN => n14427);
   U12925 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_14_7_port, B1 => 
                           n13808, B2 => REGISTERS_38_7_port, C1 => n13889, C2 
                           => REGISTERS_39_7_port, ZN => n14428);
   U12926 : OAI221_X1 port map( B1 => n10918, B2 => n13810, C1 => n10854, C2 =>
                           n13890, A => n14429, ZN => n14426);
   U12927 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_7_port, B1 => 
                           n341, B2 => REGISTERS_9_7_port, C1 => n13812, C2 => 
                           REGISTERS_16_7_port, ZN => n14429);
   U12928 : OAI221_X1 port map( B1 => n10758, B2 => n303, C1 => n10694, C2 => 
                           n13893, A => n14430, ZN => n14425);
   U12929 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_7_port, B1 => 
                           n352, B2 => REGISTERS_4_7_port, C1 => n13818, C2 => 
                           REGISTERS_11_7_port, ZN => n14430);
   U12930 : OAI221_X1 port map( B1 => n11622, B2 => n304, C1 => n10566, C2 => 
                           n13896, A => n14431, ZN => n14424);
   U12931 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_7_port, B1 => 
                           n13826, B2 => REGISTERS_0_7_port, C1 => n13824, C2 
                           => REGISTERS_6_7_port, ZN => n14431);
   U12932 : NOR4_X1 port map( A1 => n14432, A2 => n14433, A3 => n14434, A4 => 
                           n14435, ZN => n14422);
   U12933 : OAI221_X1 port map( B1 => n11686, B2 => n369, C1 => n10950, C2 => 
                           n380, A => n14436, ZN => n14435);
   U12934 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_29_7_port, B1 => 
                           n402, B2 => REGISTERS_33_7_port, C1 => n413, C2 => 
                           REGISTERS_37_7_port, ZN => n14436);
   U12935 : OAI221_X1 port map( B1 => n11526, B2 => n424, C1 => n11654, C2 => 
                           n435, A => n14437, ZN => n14434);
   U12936 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_24_7_port, B1 => 
                           n457, B2 => REGISTERS_28_7_port, C1 => n468, C2 => 
                           REGISTERS_32_7_port, ZN => n14437);
   U12937 : OAI221_X1 port map( B1 => n11366, B2 => n479, C1 => n11494, C2 => 
                           n490, A => n14438, ZN => n14433);
   U12938 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_19_7_port, B1 => 
                           n512, B2 => REGISTERS_23_7_port, C1 => n523, C2 => 
                           REGISTERS_27_7_port, ZN => n14438);
   U12939 : OAI221_X1 port map( B1 => n11206, B2 => n534, C1 => n11334, C2 => 
                           n545, A => n14439, ZN => n14432);
   U12940 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_22_7_port, B1 => 
                           n567, B2 => REGISTERS_20_7_port, C1 => n578, C2 => 
                           REGISTERS_18_7_port, ZN => n14439);
   U12941 : NOR4_X1 port map( A1 => n14442, A2 => n14443, A3 => n14444, A4 => 
                           n14445, ZN => n14441);
   U12942 : OAI221_X1 port map( B1 => n11046, B2 => n314, C1 => n10982, C2 => 
                           n325, A => n14446, ZN => n14445);
   U12943 : AOI222_X1 port map( A1 => n336, A2 => REGISTERS_13_7_port, B1 => 
                           n13808, B2 => REGISTERS_37_7_port, C1 => n13889, C2 
                           => REGISTERS_38_7_port, ZN => n14446);
   U12944 : OAI221_X1 port map( B1 => n10886, B2 => n13810, C1 => n10822, C2 =>
                           n13890, A => n14447, ZN => n14444);
   U12945 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_7_port, B1 => 
                           n343, B2 => REGISTERS_8_7_port, C1 => n13812, C2 => 
                           REGISTERS_15_7_port, ZN => n14447);
   U12946 : OAI221_X1 port map( B1 => n10726, B2 => n303, C1 => n10662, C2 => 
                           n13893, A => n14448, ZN => n14443);
   U12947 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_7_port, B1 => 
                           n354, B2 => REGISTERS_3_7_port, C1 => n13818, C2 => 
                           REGISTERS_10_7_port, ZN => n14448);
   U12948 : OAI221_X1 port map( B1 => n11590, B2 => n304, C1 => n10520, C2 => 
                           n13896, A => n14449, ZN => n14442);
   U12949 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_7_port, B1 => 
                           n13917, B2 => REGISTERS_39_7_port, C1 => n13824, C2 
                           => REGISTERS_5_7_port, ZN => n14449);
   U12950 : NOR4_X1 port map( A1 => n14450, A2 => n14451, A3 => n14452, A4 => 
                           n14453, ZN => n14440);
   U12951 : OAI221_X1 port map( B1 => n11654, B2 => n369, C1 => n10918, C2 => 
                           n380, A => n14454, ZN => n14453);
   U12952 : AOI222_X1 port map( A1 => n391, A2 => REGISTERS_28_7_port, B1 => 
                           n402, B2 => REGISTERS_32_7_port, C1 => n413, C2 => 
                           REGISTERS_36_7_port, ZN => n14454);
   U12953 : OAI221_X1 port map( B1 => n11494, B2 => n424, C1 => n11622, C2 => 
                           n435, A => n14455, ZN => n14452);
   U12954 : AOI222_X1 port map( A1 => n446, A2 => REGISTERS_23_7_port, B1 => 
                           n457, B2 => REGISTERS_27_7_port, C1 => n468, C2 => 
                           REGISTERS_31_7_port, ZN => n14455);
   U12955 : OAI221_X1 port map( B1 => n11334, B2 => n479, C1 => n11462, C2 => 
                           n490, A => n14456, ZN => n14451);
   U12956 : AOI222_X1 port map( A1 => n501, A2 => REGISTERS_18_7_port, B1 => 
                           n512, B2 => REGISTERS_22_7_port, C1 => n523, C2 => 
                           REGISTERS_26_7_port, ZN => n14456);
   U12957 : OAI221_X1 port map( B1 => n11174, B2 => n534, C1 => n11302, C2 => 
                           n545, A => n14457, ZN => n14450);
   U12958 : AOI222_X1 port map( A1 => n556, A2 => REGISTERS_21_7_port, B1 => 
                           n567, B2 => REGISTERS_19_7_port, C1 => n578, C2 => 
                           REGISTERS_17_7_port, ZN => n14457);
   U12959 : NAND3_X1 port map( A1 => n14458, A2 => n14459, A3 => n14460, ZN => 
                           n11896);
   U12960 : AOI221_X1 port map( B1 => n13792, B2 => n4949, C1 => n13793, C2 => 
                           MEM_IN(8), A => n14461, ZN => n14460);
   U12961 : OAI22_X1 port map( A1 => n10517, A2 => n251, B1 => n4951, B2 => 
                           n121, ZN => n14461);
   U12962 : NOR2_X1 port map( A1 => n5592, A2 => n13796, ZN => n5590);
   U12963 : INV_X1 port map( A => MEM_IN(8), ZN => n5592);
   U12964 : AOI22_X1 port map( A1 => n197, A2 => n4952, B1 => n150, B2 => n4953
                           , ZN => n14459);
   U12965 : NOR4_X1 port map( A1 => n14464, A2 => n14465, A3 => n14466, A4 => 
                           n14467, ZN => n14463);
   U12966 : OAI221_X1 port map( B1 => n11109, B2 => n313, C1 => n11045, C2 => 
                           n324, A => n14468, ZN => n14467);
   U12967 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_15_8_port, B1 => 
                           n13807, B2 => REGISTERS_11_8_port, C1 => n13808, C2 
                           => REGISTERS_39_8_port, ZN => n14468);
   U12968 : OAI221_X1 port map( B1 => n10821, B2 => n13809, C1 => n10949, C2 =>
                           n13810, A => n14469, ZN => n14466);
   U12969 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_8_port, B1 => 
                           n13813, B2 => REGISTERS_6_8_port, C1 => n347, C2 => 
                           REGISTERS_10_8_port, ZN => n14469);
   U12970 : OAI221_X1 port map( B1 => n10661, B2 => n13815, C1 => n10789, C2 =>
                           n303, A => n14470, ZN => n14465);
   U12971 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_8_port, B1 => 
                           n13819, B2 => REGISTERS_2_8_port, C1 => n358, C2 => 
                           REGISTERS_5_8_port, ZN => n14470);
   U12972 : OAI221_X1 port map( B1 => n10629, B2 => n13821, C1 => n11653, C2 =>
                           n304, A => n14471, ZN => n14464);
   U12973 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_8_port, B1 => 
                           n13825, B2 => REGISTERS_0_8_port, C1 => n13826, C2 
                           => REGISTERS_1_8_port, ZN => n14471);
   U12974 : NOR4_X1 port map( A1 => n14472, A2 => n14473, A3 => n14474, A4 => 
                           n14475, ZN => n14462);
   U12975 : OAI221_X1 port map( B1 => n11717, B2 => n368, C1 => n10981, C2 => 
                           n380, A => n14476, ZN => n14475);
   U12976 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_30_8_port, B1 => 
                           n401, B2 => REGISTERS_34_8_port, C1 => n412, C2 => 
                           REGISTERS_38_8_port, ZN => n14476);
   U12977 : OAI221_X1 port map( B1 => n11557, B2 => n423, C1 => n11685, C2 => 
                           n434, A => n14477, ZN => n14474);
   U12978 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_25_8_port, B1 => 
                           n456, B2 => REGISTERS_29_8_port, C1 => n467, C2 => 
                           REGISTERS_33_8_port, ZN => n14477);
   U12979 : OAI221_X1 port map( B1 => n11397, B2 => n478, C1 => n11525, C2 => 
                           n489, A => n14478, ZN => n14473);
   U12980 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_20_8_port, B1 => 
                           n511, B2 => REGISTERS_24_8_port, C1 => n522, C2 => 
                           REGISTERS_28_8_port, ZN => n14478);
   U12981 : OAI221_X1 port map( B1 => n11237, B2 => n533, C1 => n11365, C2 => 
                           n544, A => n14479, ZN => n14472);
   U12982 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_23_8_port, B1 => 
                           n566, B2 => REGISTERS_21_8_port, C1 => n577, C2 => 
                           REGISTERS_19_8_port, ZN => n14479);
   U12983 : NOR4_X1 port map( A1 => n14482, A2 => n14483, A3 => n14484, A4 => 
                           n14485, ZN => n14481);
   U12984 : OAI221_X1 port map( B1 => n11141, B2 => n313, C1 => n11077, C2 => 
                           n324, A => n14486, ZN => n14485);
   U12985 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_16_8_port, B1 => 
                           n119, B2 => REGISTERS_14_8_port, C1 => n13807, C2 =>
                           REGISTERS_12_8_port, ZN => n14486);
   U12986 : OAI221_X1 port map( B1 => n11109, B2 => n13863, C1 => n10853, C2 =>
                           n13809, A => n14487, ZN => n14484);
   U12987 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_8_port, B1 => 
                           n13865, B2 => REGISTERS_9_8_port, C1 => n13813, C2 
                           => REGISTERS_7_8_port, ZN => n14487);
   U12988 : OAI221_X1 port map( B1 => n10949, B2 => n13866, C1 => n10693, C2 =>
                           n13815, A => n14488, ZN => n14483);
   U12989 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_8_port, B1 => 
                           n13868, B2 => REGISTERS_36_8_port, C1 => n13819, C2 
                           => REGISTERS_3_8_port, ZN => n14488);
   U12990 : OAI221_X1 port map( B1 => n10789, B2 => n13869, C1 => n10661, C2 =>
                           n13821, A => n14489, ZN => n14482);
   U12991 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_8_port, B1 => 
                           n13871, B2 => REGISTERS_0_8_port, C1 => n13825, C2 
                           => REGISTERS_1_8_port, ZN => n14489);
   U12992 : NOR4_X1 port map( A1 => n14490, A2 => n14491, A3 => n14492, A4 => 
                           n14493, ZN => n14480);
   U12993 : OAI221_X1 port map( B1 => n11749, B2 => n368, C1 => n11013, C2 => 
                           n379, A => n14494, ZN => n14493);
   U12994 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_31_8_port, B1 => 
                           n401, B2 => REGISTERS_35_8_port, C1 => n412, C2 => 
                           REGISTERS_39_8_port, ZN => n14494);
   U12995 : OAI221_X1 port map( B1 => n11589, B2 => n423, C1 => n11717, C2 => 
                           n434, A => n14495, ZN => n14492);
   U12996 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_26_8_port, B1 => 
                           n456, B2 => REGISTERS_30_8_port, C1 => n467, C2 => 
                           REGISTERS_34_8_port, ZN => n14495);
   U12997 : OAI221_X1 port map( B1 => n11429, B2 => n478, C1 => n11557, C2 => 
                           n489, A => n14496, ZN => n14491);
   U12998 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_21_8_port, B1 => 
                           n511, B2 => REGISTERS_25_8_port, C1 => n522, C2 => 
                           REGISTERS_29_8_port, ZN => n14496);
   U12999 : OAI221_X1 port map( B1 => n11269, B2 => n533, C1 => n11397, C2 => 
                           n544, A => n14497, ZN => n14490);
   U13000 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_24_8_port, B1 => 
                           n566, B2 => REGISTERS_22_8_port, C1 => n577, C2 => 
                           REGISTERS_20_8_port, ZN => n14497);
   U13001 : AOI22_X1 port map( A1 => n13880, A2 => n4954, B1 => n13881, B2 => 
                           n4955, ZN => n14458);
   U13002 : NOR4_X1 port map( A1 => n14500, A2 => n14501, A3 => n14502, A4 => 
                           n14503, ZN => n14499);
   U13003 : OAI221_X1 port map( B1 => n11077, B2 => n313, C1 => n11013, C2 => 
                           n324, A => n14504, ZN => n14503);
   U13004 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_14_8_port, B1 => 
                           n13808, B2 => REGISTERS_38_8_port, C1 => n13889, C2 
                           => REGISTERS_39_8_port, ZN => n14504);
   U13005 : OAI221_X1 port map( B1 => n10917, B2 => n13810, C1 => n10853, C2 =>
                           n13890, A => n14505, ZN => n14502);
   U13006 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_8_port, B1 => 
                           n342, B2 => REGISTERS_9_8_port, C1 => n13812, C2 => 
                           REGISTERS_16_8_port, ZN => n14505);
   U13007 : OAI221_X1 port map( B1 => n10757, B2 => n303, C1 => n10693, C2 => 
                           n13893, A => n14506, ZN => n14501);
   U13008 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_8_port, B1 => 
                           n353, B2 => REGISTERS_4_8_port, C1 => n13818, C2 => 
                           REGISTERS_11_8_port, ZN => n14506);
   U13009 : OAI221_X1 port map( B1 => n11621, B2 => n304, C1 => n10565, C2 => 
                           n13896, A => n14507, ZN => n14500);
   U13010 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_8_port, B1 => 
                           n13826, B2 => REGISTERS_0_8_port, C1 => n13824, C2 
                           => REGISTERS_6_8_port, ZN => n14507);
   U13011 : NOR4_X1 port map( A1 => n14508, A2 => n14509, A3 => n14510, A4 => 
                           n14511, ZN => n14498);
   U13012 : OAI221_X1 port map( B1 => n11685, B2 => n368, C1 => n10949, C2 => 
                           n379, A => n14512, ZN => n14511);
   U13013 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_29_8_port, B1 => 
                           n401, B2 => REGISTERS_33_8_port, C1 => n412, C2 => 
                           REGISTERS_37_8_port, ZN => n14512);
   U13014 : OAI221_X1 port map( B1 => n11525, B2 => n423, C1 => n11653, C2 => 
                           n434, A => n14513, ZN => n14510);
   U13015 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_24_8_port, B1 => 
                           n456, B2 => REGISTERS_28_8_port, C1 => n467, C2 => 
                           REGISTERS_32_8_port, ZN => n14513);
   U13016 : OAI221_X1 port map( B1 => n11365, B2 => n478, C1 => n11493, C2 => 
                           n489, A => n14514, ZN => n14509);
   U13017 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_19_8_port, B1 => 
                           n511, B2 => REGISTERS_23_8_port, C1 => n522, C2 => 
                           REGISTERS_27_8_port, ZN => n14514);
   U13018 : OAI221_X1 port map( B1 => n11205, B2 => n533, C1 => n11333, C2 => 
                           n544, A => n14515, ZN => n14508);
   U13019 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_22_8_port, B1 => 
                           n566, B2 => REGISTERS_20_8_port, C1 => n577, C2 => 
                           REGISTERS_18_8_port, ZN => n14515);
   U13020 : NOR4_X1 port map( A1 => n14518, A2 => n14519, A3 => n14520, A4 => 
                           n14521, ZN => n14517);
   U13021 : OAI221_X1 port map( B1 => n11045, B2 => n313, C1 => n10981, C2 => 
                           n324, A => n14522, ZN => n14521);
   U13022 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_13_8_port, B1 => 
                           n13808, B2 => REGISTERS_37_8_port, C1 => n13889, C2 
                           => REGISTERS_38_8_port, ZN => n14522);
   U13023 : OAI221_X1 port map( B1 => n10885, B2 => n13810, C1 => n10821, C2 =>
                           n13890, A => n14523, ZN => n14520);
   U13024 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_8_port, B1 => 
                           n342, B2 => REGISTERS_8_8_port, C1 => n13812, C2 => 
                           REGISTERS_15_8_port, ZN => n14523);
   U13025 : OAI221_X1 port map( B1 => n10725, B2 => n303, C1 => n10661, C2 => 
                           n13893, A => n14524, ZN => n14519);
   U13026 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_8_port, B1 => 
                           n353, B2 => REGISTERS_3_8_port, C1 => n13818, C2 => 
                           REGISTERS_10_8_port, ZN => n14524);
   U13027 : OAI221_X1 port map( B1 => n11589, B2 => n304, C1 => n10517, C2 => 
                           n13896, A => n14525, ZN => n14518);
   U13028 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_8_port, B1 => 
                           n13917, B2 => REGISTERS_39_8_port, C1 => n13824, C2 
                           => REGISTERS_5_8_port, ZN => n14525);
   U13029 : NOR4_X1 port map( A1 => n14526, A2 => n14527, A3 => n14528, A4 => 
                           n14529, ZN => n14516);
   U13030 : OAI221_X1 port map( B1 => n11653, B2 => n368, C1 => n10917, C2 => 
                           n379, A => n14530, ZN => n14529);
   U13031 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_28_8_port, B1 => 
                           n401, B2 => REGISTERS_32_8_port, C1 => n412, C2 => 
                           REGISTERS_36_8_port, ZN => n14530);
   U13032 : OAI221_X1 port map( B1 => n11493, B2 => n423, C1 => n11621, C2 => 
                           n434, A => n14531, ZN => n14528);
   U13033 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_23_8_port, B1 => 
                           n456, B2 => REGISTERS_27_8_port, C1 => n467, C2 => 
                           REGISTERS_31_8_port, ZN => n14531);
   U13034 : OAI221_X1 port map( B1 => n11333, B2 => n478, C1 => n11461, C2 => 
                           n489, A => n14532, ZN => n14527);
   U13035 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_18_8_port, B1 => 
                           n511, B2 => REGISTERS_22_8_port, C1 => n522, C2 => 
                           REGISTERS_26_8_port, ZN => n14532);
   U13036 : OAI221_X1 port map( B1 => n11173, B2 => n533, C1 => n11301, C2 => 
                           n544, A => n14533, ZN => n14526);
   U13037 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_21_8_port, B1 => 
                           n566, B2 => REGISTERS_19_8_port, C1 => n577, C2 => 
                           REGISTERS_17_8_port, ZN => n14533);
   U13038 : NAND3_X1 port map( A1 => n14534, A2 => n14535, A3 => n14536, ZN => 
                           n11895);
   U13039 : AOI221_X1 port map( B1 => n13792, B2 => n4959, C1 => n13793, C2 => 
                           MEM_IN(9), A => n14537, ZN => n14536);
   U13040 : OAI22_X1 port map( A1 => n10514, A2 => n251, B1 => n4961, B2 => 
                           n121, ZN => n14537);
   U13041 : NOR2_X1 port map( A1 => n5599, A2 => n13796, ZN => n5597);
   U13042 : INV_X1 port map( A => MEM_IN(9), ZN => n5599);
   U13043 : AOI22_X1 port map( A1 => n197, A2 => n4962, B1 => n150, B2 => n4963
                           , ZN => n14535);
   U13044 : NOR4_X1 port map( A1 => n14540, A2 => n14541, A3 => n14542, A4 => 
                           n14543, ZN => n14539);
   U13045 : OAI221_X1 port map( B1 => n11108, B2 => n313, C1 => n11044, C2 => 
                           n324, A => n14544, ZN => n14543);
   U13046 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_15_9_port, B1 => 
                           n13807, B2 => REGISTERS_11_9_port, C1 => n13808, C2 
                           => REGISTERS_39_9_port, ZN => n14544);
   U13047 : OAI221_X1 port map( B1 => n10820, B2 => n13809, C1 => n10948, C2 =>
                           n13810, A => n14545, ZN => n14542);
   U13048 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_9_port, B1 => 
                           n13813, B2 => REGISTERS_6_9_port, C1 => n347, C2 => 
                           REGISTERS_10_9_port, ZN => n14545);
   U13049 : OAI221_X1 port map( B1 => n10660, B2 => n13815, C1 => n10788, C2 =>
                           n303, A => n14546, ZN => n14541);
   U13050 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_9_port, B1 => 
                           n13819, B2 => REGISTERS_2_9_port, C1 => n358, C2 => 
                           REGISTERS_5_9_port, ZN => n14546);
   U13051 : OAI221_X1 port map( B1 => n10628, B2 => n13821, C1 => n11652, C2 =>
                           n304, A => n14547, ZN => n14540);
   U13052 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_9_port, B1 => 
                           n13825, B2 => REGISTERS_0_9_port, C1 => n13826, C2 
                           => REGISTERS_1_9_port, ZN => n14547);
   U13053 : NOR4_X1 port map( A1 => n14548, A2 => n14549, A3 => n14550, A4 => 
                           n14551, ZN => n14538);
   U13054 : OAI221_X1 port map( B1 => n11716, B2 => n368, C1 => n10980, C2 => 
                           n379, A => n14552, ZN => n14551);
   U13055 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_30_9_port, B1 => 
                           n401, B2 => REGISTERS_34_9_port, C1 => n412, C2 => 
                           REGISTERS_38_9_port, ZN => n14552);
   U13056 : OAI221_X1 port map( B1 => n11556, B2 => n423, C1 => n11684, C2 => 
                           n434, A => n14553, ZN => n14550);
   U13057 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_25_9_port, B1 => 
                           n456, B2 => REGISTERS_29_9_port, C1 => n467, C2 => 
                           REGISTERS_33_9_port, ZN => n14553);
   U13058 : OAI221_X1 port map( B1 => n11396, B2 => n478, C1 => n11524, C2 => 
                           n489, A => n14554, ZN => n14549);
   U13059 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_20_9_port, B1 => 
                           n511, B2 => REGISTERS_24_9_port, C1 => n522, C2 => 
                           REGISTERS_28_9_port, ZN => n14554);
   U13060 : OAI221_X1 port map( B1 => n11236, B2 => n533, C1 => n11364, C2 => 
                           n544, A => n14555, ZN => n14548);
   U13061 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_23_9_port, B1 => 
                           n566, B2 => REGISTERS_21_9_port, C1 => n577, C2 => 
                           REGISTERS_19_9_port, ZN => n14555);
   U13062 : NOR4_X1 port map( A1 => n14558, A2 => n14559, A3 => n14560, A4 => 
                           n14561, ZN => n14557);
   U13063 : OAI221_X1 port map( B1 => n11140, B2 => n313, C1 => n11076, C2 => 
                           n324, A => n14562, ZN => n14561);
   U13064 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_16_9_port, B1 => 
                           n119, B2 => REGISTERS_14_9_port, C1 => n13807, C2 =>
                           REGISTERS_12_9_port, ZN => n14562);
   U13065 : OAI221_X1 port map( B1 => n11108, B2 => n13863, C1 => n10852, C2 =>
                           n13809, A => n14563, ZN => n14560);
   U13066 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_9_port, B1 => 
                           n13865, B2 => REGISTERS_9_9_port, C1 => n13813, C2 
                           => REGISTERS_7_9_port, ZN => n14563);
   U13067 : OAI221_X1 port map( B1 => n10948, B2 => n13866, C1 => n10692, C2 =>
                           n13815, A => n14564, ZN => n14559);
   U13068 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_9_port, B1 => 
                           n13868, B2 => REGISTERS_36_9_port, C1 => n13819, C2 
                           => REGISTERS_3_9_port, ZN => n14564);
   U13069 : OAI221_X1 port map( B1 => n10788, B2 => n13869, C1 => n10660, C2 =>
                           n13821, A => n14565, ZN => n14558);
   U13070 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_9_port, B1 => 
                           n13871, B2 => REGISTERS_0_9_port, C1 => n13825, C2 
                           => REGISTERS_1_9_port, ZN => n14565);
   U13071 : NOR4_X1 port map( A1 => n14566, A2 => n14567, A3 => n14568, A4 => 
                           n14569, ZN => n14556);
   U13072 : OAI221_X1 port map( B1 => n11748, B2 => n368, C1 => n11012, C2 => 
                           n379, A => n14570, ZN => n14569);
   U13073 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_31_9_port, B1 => 
                           n401, B2 => REGISTERS_35_9_port, C1 => n412, C2 => 
                           REGISTERS_39_9_port, ZN => n14570);
   U13074 : OAI221_X1 port map( B1 => n11588, B2 => n423, C1 => n11716, C2 => 
                           n434, A => n14571, ZN => n14568);
   U13075 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_26_9_port, B1 => 
                           n456, B2 => REGISTERS_30_9_port, C1 => n467, C2 => 
                           REGISTERS_34_9_port, ZN => n14571);
   U13076 : OAI221_X1 port map( B1 => n11428, B2 => n478, C1 => n11556, C2 => 
                           n489, A => n14572, ZN => n14567);
   U13077 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_21_9_port, B1 => 
                           n511, B2 => REGISTERS_25_9_port, C1 => n522, C2 => 
                           REGISTERS_29_9_port, ZN => n14572);
   U13078 : OAI221_X1 port map( B1 => n11268, B2 => n533, C1 => n11396, C2 => 
                           n544, A => n14573, ZN => n14566);
   U13079 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_24_9_port, B1 => 
                           n566, B2 => REGISTERS_22_9_port, C1 => n577, C2 => 
                           REGISTERS_20_9_port, ZN => n14573);
   U13080 : AOI22_X1 port map( A1 => n13880, A2 => n4964, B1 => n13881, B2 => 
                           n4965, ZN => n14534);
   U13081 : NOR4_X1 port map( A1 => n14576, A2 => n14577, A3 => n14578, A4 => 
                           n14579, ZN => n14575);
   U13082 : OAI221_X1 port map( B1 => n11076, B2 => n313, C1 => n11012, C2 => 
                           n324, A => n14580, ZN => n14579);
   U13083 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_14_9_port, B1 => 
                           n13808, B2 => REGISTERS_38_9_port, C1 => n13889, C2 
                           => REGISTERS_39_9_port, ZN => n14580);
   U13084 : OAI221_X1 port map( B1 => n10916, B2 => n13810, C1 => n10852, C2 =>
                           n13890, A => n14581, ZN => n14578);
   U13085 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_9_port, B1 => 
                           n343, B2 => REGISTERS_9_9_port, C1 => n13812, C2 => 
                           REGISTERS_16_9_port, ZN => n14581);
   U13086 : OAI221_X1 port map( B1 => n10756, B2 => n303, C1 => n10692, C2 => 
                           n13893, A => n14582, ZN => n14577);
   U13087 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_9_port, B1 => 
                           n354, B2 => REGISTERS_4_9_port, C1 => n13818, C2 => 
                           REGISTERS_11_9_port, ZN => n14582);
   U13088 : OAI221_X1 port map( B1 => n11620, B2 => n304, C1 => n10564, C2 => 
                           n13896, A => n14583, ZN => n14576);
   U13089 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_9_port, B1 => 
                           n13826, B2 => REGISTERS_0_9_port, C1 => n13824, C2 
                           => REGISTERS_6_9_port, ZN => n14583);
   U13090 : NOR4_X1 port map( A1 => n14584, A2 => n14585, A3 => n14586, A4 => 
                           n14587, ZN => n14574);
   U13091 : OAI221_X1 port map( B1 => n11684, B2 => n368, C1 => n10948, C2 => 
                           n379, A => n14588, ZN => n14587);
   U13092 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_29_9_port, B1 => 
                           n401, B2 => REGISTERS_33_9_port, C1 => n412, C2 => 
                           REGISTERS_37_9_port, ZN => n14588);
   U13093 : OAI221_X1 port map( B1 => n11524, B2 => n423, C1 => n11652, C2 => 
                           n434, A => n14589, ZN => n14586);
   U13094 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_24_9_port, B1 => 
                           n456, B2 => REGISTERS_28_9_port, C1 => n467, C2 => 
                           REGISTERS_32_9_port, ZN => n14589);
   U13095 : OAI221_X1 port map( B1 => n11364, B2 => n478, C1 => n11492, C2 => 
                           n489, A => n14590, ZN => n14585);
   U13096 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_19_9_port, B1 => 
                           n511, B2 => REGISTERS_23_9_port, C1 => n522, C2 => 
                           REGISTERS_27_9_port, ZN => n14590);
   U13097 : OAI221_X1 port map( B1 => n11204, B2 => n533, C1 => n11332, C2 => 
                           n544, A => n14591, ZN => n14584);
   U13098 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_22_9_port, B1 => 
                           n566, B2 => REGISTERS_20_9_port, C1 => n577, C2 => 
                           REGISTERS_18_9_port, ZN => n14591);
   U13099 : NOR4_X1 port map( A1 => n14594, A2 => n14595, A3 => n14596, A4 => 
                           n14597, ZN => n14593);
   U13100 : OAI221_X1 port map( B1 => n11044, B2 => n313, C1 => n10980, C2 => 
                           n324, A => n14598, ZN => n14597);
   U13101 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_13_9_port, B1 => 
                           n13808, B2 => REGISTERS_37_9_port, C1 => n13889, C2 
                           => REGISTERS_38_9_port, ZN => n14598);
   U13102 : OAI221_X1 port map( B1 => n10884, B2 => n13810, C1 => n10820, C2 =>
                           n13890, A => n14599, ZN => n14596);
   U13103 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_9_port, B1 => 
                           n341, B2 => REGISTERS_8_9_port, C1 => n13812, C2 => 
                           REGISTERS_15_9_port, ZN => n14599);
   U13104 : OAI221_X1 port map( B1 => n10724, B2 => n303, C1 => n10660, C2 => 
                           n13893, A => n14600, ZN => n14595);
   U13105 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_9_port, B1 => 
                           n352, B2 => REGISTERS_3_9_port, C1 => n13818, C2 => 
                           REGISTERS_10_9_port, ZN => n14600);
   U13106 : OAI221_X1 port map( B1 => n11588, B2 => n304, C1 => n10514, C2 => 
                           n13896, A => n14601, ZN => n14594);
   U13107 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_9_port, B1 => 
                           n13917, B2 => REGISTERS_39_9_port, C1 => n13824, C2 
                           => REGISTERS_5_9_port, ZN => n14601);
   U13108 : NOR4_X1 port map( A1 => n14602, A2 => n14603, A3 => n14604, A4 => 
                           n14605, ZN => n14592);
   U13109 : OAI221_X1 port map( B1 => n11652, B2 => n368, C1 => n10916, C2 => 
                           n379, A => n14606, ZN => n14605);
   U13110 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_28_9_port, B1 => 
                           n401, B2 => REGISTERS_32_9_port, C1 => n412, C2 => 
                           REGISTERS_36_9_port, ZN => n14606);
   U13111 : OAI221_X1 port map( B1 => n11492, B2 => n423, C1 => n11620, C2 => 
                           n434, A => n14607, ZN => n14604);
   U13112 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_23_9_port, B1 => 
                           n456, B2 => REGISTERS_27_9_port, C1 => n467, C2 => 
                           REGISTERS_31_9_port, ZN => n14607);
   U13113 : OAI221_X1 port map( B1 => n11332, B2 => n478, C1 => n11460, C2 => 
                           n489, A => n14608, ZN => n14603);
   U13114 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_18_9_port, B1 => 
                           n511, B2 => REGISTERS_22_9_port, C1 => n522, C2 => 
                           REGISTERS_26_9_port, ZN => n14608);
   U13115 : OAI221_X1 port map( B1 => n11172, B2 => n533, C1 => n11300, C2 => 
                           n544, A => n14609, ZN => n14602);
   U13116 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_21_9_port, B1 => 
                           n566, B2 => REGISTERS_19_9_port, C1 => n577, C2 => 
                           REGISTERS_17_9_port, ZN => n14609);
   U13117 : NAND3_X1 port map( A1 => n14610, A2 => n14611, A3 => n14612, ZN => 
                           n11894);
   U13118 : AOI221_X1 port map( B1 => n13792, B2 => n4969, C1 => n13793, C2 => 
                           MEM_IN(10), A => n14613, ZN => n14612);
   U13119 : OAI22_X1 port map( A1 => n10511, A2 => n251, B1 => n4971, B2 => 
                           n121, ZN => n14613);
   U13120 : NOR2_X1 port map( A1 => n5606, A2 => n13796, ZN => n5604);
   U13121 : INV_X1 port map( A => MEM_IN(10), ZN => n5606);
   U13122 : AOI22_X1 port map( A1 => n197, A2 => n4972, B1 => n150, B2 => n4973
                           , ZN => n14611);
   U13123 : NOR4_X1 port map( A1 => n14616, A2 => n14617, A3 => n14618, A4 => 
                           n14619, ZN => n14615);
   U13124 : OAI221_X1 port map( B1 => n11107, B2 => n313, C1 => n11043, C2 => 
                           n324, A => n14620, ZN => n14619);
   U13125 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_15_10_port, B1 => 
                           n13807, B2 => REGISTERS_11_10_port, C1 => n13808, C2
                           => REGISTERS_39_10_port, ZN => n14620);
   U13126 : OAI221_X1 port map( B1 => n10819, B2 => n13809, C1 => n10947, C2 =>
                           n13810, A => n14621, ZN => n14618);
   U13127 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_10_port, B1 =>
                           n13813, B2 => REGISTERS_6_10_port, C1 => n347, C2 =>
                           REGISTERS_10_10_port, ZN => n14621);
   U13128 : OAI221_X1 port map( B1 => n10659, B2 => n13815, C1 => n10787, C2 =>
                           n303, A => n14622, ZN => n14617);
   U13129 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_10_port, B1 =>
                           n13819, B2 => REGISTERS_2_10_port, C1 => n358, C2 =>
                           REGISTERS_5_10_port, ZN => n14622);
   U13130 : OAI221_X1 port map( B1 => n10627, B2 => n13821, C1 => n11651, C2 =>
                           n304, A => n14623, ZN => n14616);
   U13131 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_10_port, B1 => 
                           n13825, B2 => REGISTERS_0_10_port, C1 => n13826, C2 
                           => REGISTERS_1_10_port, ZN => n14623);
   U13132 : NOR4_X1 port map( A1 => n14624, A2 => n14625, A3 => n14626, A4 => 
                           n14627, ZN => n14614);
   U13133 : OAI221_X1 port map( B1 => n11715, B2 => n368, C1 => n10979, C2 => 
                           n379, A => n14628, ZN => n14627);
   U13134 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_30_10_port, B1 => 
                           n401, B2 => REGISTERS_34_10_port, C1 => n412, C2 => 
                           REGISTERS_38_10_port, ZN => n14628);
   U13135 : OAI221_X1 port map( B1 => n11555, B2 => n423, C1 => n11683, C2 => 
                           n434, A => n14629, ZN => n14626);
   U13136 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_25_10_port, B1 => 
                           n456, B2 => REGISTERS_29_10_port, C1 => n467, C2 => 
                           REGISTERS_33_10_port, ZN => n14629);
   U13137 : OAI221_X1 port map( B1 => n11395, B2 => n478, C1 => n11523, C2 => 
                           n489, A => n14630, ZN => n14625);
   U13138 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_20_10_port, B1 => 
                           n511, B2 => REGISTERS_24_10_port, C1 => n522, C2 => 
                           REGISTERS_28_10_port, ZN => n14630);
   U13139 : OAI221_X1 port map( B1 => n11235, B2 => n533, C1 => n11363, C2 => 
                           n544, A => n14631, ZN => n14624);
   U13140 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_23_10_port, B1 => 
                           n566, B2 => REGISTERS_21_10_port, C1 => n577, C2 => 
                           REGISTERS_19_10_port, ZN => n14631);
   U13141 : NOR4_X1 port map( A1 => n14634, A2 => n14635, A3 => n14636, A4 => 
                           n14637, ZN => n14633);
   U13142 : OAI221_X1 port map( B1 => n11139, B2 => n313, C1 => n11075, C2 => 
                           n324, A => n14638, ZN => n14637);
   U13143 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_16_10_port, B1 => 
                           n119, B2 => REGISTERS_14_10_port, C1 => n13807, C2 
                           => REGISTERS_12_10_port, ZN => n14638);
   U13144 : OAI221_X1 port map( B1 => n11107, B2 => n13863, C1 => n10851, C2 =>
                           n13809, A => n14639, ZN => n14636);
   U13145 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_10_port, B1 => 
                           n13865, B2 => REGISTERS_9_10_port, C1 => n13813, C2 
                           => REGISTERS_7_10_port, ZN => n14639);
   U13146 : OAI221_X1 port map( B1 => n10947, B2 => n13866, C1 => n10691, C2 =>
                           n13815, A => n14640, ZN => n14635);
   U13147 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_10_port, B1 => 
                           n13868, B2 => REGISTERS_36_10_port, C1 => n13819, C2
                           => REGISTERS_3_10_port, ZN => n14640);
   U13148 : OAI221_X1 port map( B1 => n10787, B2 => n13869, C1 => n10659, C2 =>
                           n13821, A => n14641, ZN => n14634);
   U13149 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_10_port, B1 => 
                           n13871, B2 => REGISTERS_0_10_port, C1 => n13825, C2 
                           => REGISTERS_1_10_port, ZN => n14641);
   U13150 : NOR4_X1 port map( A1 => n14642, A2 => n14643, A3 => n14644, A4 => 
                           n14645, ZN => n14632);
   U13151 : OAI221_X1 port map( B1 => n11747, B2 => n368, C1 => n11011, C2 => 
                           n379, A => n14646, ZN => n14645);
   U13152 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_31_10_port, B1 => 
                           n401, B2 => REGISTERS_35_10_port, C1 => n412, C2 => 
                           REGISTERS_39_10_port, ZN => n14646);
   U13153 : OAI221_X1 port map( B1 => n11587, B2 => n423, C1 => n11715, C2 => 
                           n434, A => n14647, ZN => n14644);
   U13154 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_26_10_port, B1 => 
                           n456, B2 => REGISTERS_30_10_port, C1 => n467, C2 => 
                           REGISTERS_34_10_port, ZN => n14647);
   U13155 : OAI221_X1 port map( B1 => n11427, B2 => n478, C1 => n11555, C2 => 
                           n489, A => n14648, ZN => n14643);
   U13156 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_21_10_port, B1 => 
                           n511, B2 => REGISTERS_25_10_port, C1 => n522, C2 => 
                           REGISTERS_29_10_port, ZN => n14648);
   U13157 : OAI221_X1 port map( B1 => n11267, B2 => n533, C1 => n11395, C2 => 
                           n544, A => n14649, ZN => n14642);
   U13158 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_24_10_port, B1 => 
                           n566, B2 => REGISTERS_22_10_port, C1 => n577, C2 => 
                           REGISTERS_20_10_port, ZN => n14649);
   U13159 : AOI22_X1 port map( A1 => n13880, A2 => n4974, B1 => n13881, B2 => 
                           n4975, ZN => n14610);
   U13160 : NOR4_X1 port map( A1 => n14652, A2 => n14653, A3 => n14654, A4 => 
                           n14655, ZN => n14651);
   U13161 : OAI221_X1 port map( B1 => n11075, B2 => n313, C1 => n11011, C2 => 
                           n324, A => n14656, ZN => n14655);
   U13162 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_14_10_port, B1 => 
                           n13808, B2 => REGISTERS_38_10_port, C1 => n13889, C2
                           => REGISTERS_39_10_port, ZN => n14656);
   U13163 : OAI221_X1 port map( B1 => n10915, B2 => n13810, C1 => n10851, C2 =>
                           n13890, A => n14657, ZN => n14654);
   U13164 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_10_port, B1 => 
                           n342, B2 => REGISTERS_9_10_port, C1 => n13812, C2 =>
                           REGISTERS_16_10_port, ZN => n14657);
   U13165 : OAI221_X1 port map( B1 => n10755, B2 => n303, C1 => n10691, C2 => 
                           n13893, A => n14658, ZN => n14653);
   U13166 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_10_port, B1 => 
                           n353, B2 => REGISTERS_4_10_port, C1 => n13818, C2 =>
                           REGISTERS_11_10_port, ZN => n14658);
   U13167 : OAI221_X1 port map( B1 => n11619, B2 => n304, C1 => n10563, C2 => 
                           n13896, A => n14659, ZN => n14652);
   U13168 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_10_port, B1 => 
                           n13826, B2 => REGISTERS_0_10_port, C1 => n13824, C2 
                           => REGISTERS_6_10_port, ZN => n14659);
   U13169 : NOR4_X1 port map( A1 => n14660, A2 => n14661, A3 => n14662, A4 => 
                           n14663, ZN => n14650);
   U13170 : OAI221_X1 port map( B1 => n11683, B2 => n368, C1 => n10947, C2 => 
                           n379, A => n14664, ZN => n14663);
   U13171 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_29_10_port, B1 => 
                           n401, B2 => REGISTERS_33_10_port, C1 => n412, C2 => 
                           REGISTERS_37_10_port, ZN => n14664);
   U13172 : OAI221_X1 port map( B1 => n11523, B2 => n423, C1 => n11651, C2 => 
                           n434, A => n14665, ZN => n14662);
   U13173 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_24_10_port, B1 => 
                           n456, B2 => REGISTERS_28_10_port, C1 => n467, C2 => 
                           REGISTERS_32_10_port, ZN => n14665);
   U13174 : OAI221_X1 port map( B1 => n11363, B2 => n478, C1 => n11491, C2 => 
                           n489, A => n14666, ZN => n14661);
   U13175 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_19_10_port, B1 => 
                           n511, B2 => REGISTERS_23_10_port, C1 => n522, C2 => 
                           REGISTERS_27_10_port, ZN => n14666);
   U13176 : OAI221_X1 port map( B1 => n11203, B2 => n533, C1 => n11331, C2 => 
                           n544, A => n14667, ZN => n14660);
   U13177 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_22_10_port, B1 => 
                           n566, B2 => REGISTERS_20_10_port, C1 => n577, C2 => 
                           REGISTERS_18_10_port, ZN => n14667);
   U13178 : NOR4_X1 port map( A1 => n14670, A2 => n14671, A3 => n14672, A4 => 
                           n14673, ZN => n14669);
   U13179 : OAI221_X1 port map( B1 => n11043, B2 => n313, C1 => n10979, C2 => 
                           n324, A => n14674, ZN => n14673);
   U13180 : AOI222_X1 port map( A1 => n335, A2 => REGISTERS_13_10_port, B1 => 
                           n13808, B2 => REGISTERS_37_10_port, C1 => n13889, C2
                           => REGISTERS_38_10_port, ZN => n14674);
   U13181 : OAI221_X1 port map( B1 => n10883, B2 => n13810, C1 => n10819, C2 =>
                           n13890, A => n14675, ZN => n14672);
   U13182 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_10_port, B1 => 
                           n342, B2 => REGISTERS_8_10_port, C1 => n13812, C2 =>
                           REGISTERS_15_10_port, ZN => n14675);
   U13183 : OAI221_X1 port map( B1 => n10723, B2 => n303, C1 => n10659, C2 => 
                           n13893, A => n14676, ZN => n14671);
   U13184 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_10_port, B1 => 
                           n353, B2 => REGISTERS_3_10_port, C1 => n13818, C2 =>
                           REGISTERS_10_10_port, ZN => n14676);
   U13185 : OAI221_X1 port map( B1 => n11587, B2 => n304, C1 => n10511, C2 => 
                           n13896, A => n14677, ZN => n14670);
   U13186 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_10_port, B1 => 
                           n13917, B2 => REGISTERS_39_10_port, C1 => n13824, C2
                           => REGISTERS_5_10_port, ZN => n14677);
   U13187 : NOR4_X1 port map( A1 => n14678, A2 => n14679, A3 => n14680, A4 => 
                           n14681, ZN => n14668);
   U13188 : OAI221_X1 port map( B1 => n11651, B2 => n368, C1 => n10915, C2 => 
                           n379, A => n14682, ZN => n14681);
   U13189 : AOI222_X1 port map( A1 => n390, A2 => REGISTERS_28_10_port, B1 => 
                           n401, B2 => REGISTERS_32_10_port, C1 => n412, C2 => 
                           REGISTERS_36_10_port, ZN => n14682);
   U13190 : OAI221_X1 port map( B1 => n11491, B2 => n423, C1 => n11619, C2 => 
                           n434, A => n14683, ZN => n14680);
   U13191 : AOI222_X1 port map( A1 => n445, A2 => REGISTERS_23_10_port, B1 => 
                           n456, B2 => REGISTERS_27_10_port, C1 => n467, C2 => 
                           REGISTERS_31_10_port, ZN => n14683);
   U13192 : OAI221_X1 port map( B1 => n11331, B2 => n478, C1 => n11459, C2 => 
                           n489, A => n14684, ZN => n14679);
   U13193 : AOI222_X1 port map( A1 => n500, A2 => REGISTERS_18_10_port, B1 => 
                           n511, B2 => REGISTERS_22_10_port, C1 => n522, C2 => 
                           REGISTERS_26_10_port, ZN => n14684);
   U13194 : OAI221_X1 port map( B1 => n11171, B2 => n533, C1 => n11299, C2 => 
                           n544, A => n14685, ZN => n14678);
   U13195 : AOI222_X1 port map( A1 => n555, A2 => REGISTERS_21_10_port, B1 => 
                           n566, B2 => REGISTERS_19_10_port, C1 => n577, C2 => 
                           REGISTERS_17_10_port, ZN => n14685);
   U13196 : NAND3_X1 port map( A1 => n14686, A2 => n14687, A3 => n14688, ZN => 
                           n11893);
   U13197 : AOI221_X1 port map( B1 => n13792, B2 => n4979, C1 => n13793, C2 => 
                           MEM_IN(11), A => n14689, ZN => n14688);
   U13198 : OAI22_X1 port map( A1 => n10508, A2 => n251, B1 => n4981, B2 => 
                           n121, ZN => n14689);
   U13199 : NOR2_X1 port map( A1 => n5613, A2 => n13796, ZN => n5611);
   U13200 : INV_X1 port map( A => MEM_IN(11), ZN => n5613);
   U13201 : AOI22_X1 port map( A1 => n197, A2 => n4982, B1 => n150, B2 => n4983
                           , ZN => n14687);
   U13202 : NOR4_X1 port map( A1 => n14692, A2 => n14693, A3 => n14694, A4 => 
                           n14695, ZN => n14691);
   U13203 : OAI221_X1 port map( B1 => n11106, B2 => n312, C1 => n11042, C2 => 
                           n323, A => n14696, ZN => n14695);
   U13204 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_15_11_port, B1 => 
                           n13807, B2 => REGISTERS_11_11_port, C1 => n13808, C2
                           => REGISTERS_39_11_port, ZN => n14696);
   U13205 : OAI221_X1 port map( B1 => n10818, B2 => n13809, C1 => n10946, C2 =>
                           n13810, A => n14697, ZN => n14694);
   U13206 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_11_port, B1 =>
                           n13813, B2 => REGISTERS_6_11_port, C1 => n348, C2 =>
                           REGISTERS_10_11_port, ZN => n14697);
   U13207 : OAI221_X1 port map( B1 => n10658, B2 => n13815, C1 => n10786, C2 =>
                           n303, A => n14698, ZN => n14693);
   U13208 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_11_port, B1 =>
                           n13819, B2 => REGISTERS_2_11_port, C1 => n359, C2 =>
                           REGISTERS_5_11_port, ZN => n14698);
   U13209 : OAI221_X1 port map( B1 => n10626, B2 => n13821, C1 => n11650, C2 =>
                           n304, A => n14699, ZN => n14692);
   U13210 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_11_port, B1 => 
                           n13825, B2 => REGISTERS_0_11_port, C1 => n13826, C2 
                           => REGISTERS_1_11_port, ZN => n14699);
   U13211 : NOR4_X1 port map( A1 => n14700, A2 => n14701, A3 => n14702, A4 => 
                           n14703, ZN => n14690);
   U13212 : OAI221_X1 port map( B1 => n11714, B2 => n367, C1 => n10978, C2 => 
                           n379, A => n14704, ZN => n14703);
   U13213 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_30_11_port, B1 => 
                           n400, B2 => REGISTERS_34_11_port, C1 => n411, C2 => 
                           REGISTERS_38_11_port, ZN => n14704);
   U13214 : OAI221_X1 port map( B1 => n11554, B2 => n422, C1 => n11682, C2 => 
                           n433, A => n14705, ZN => n14702);
   U13215 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_25_11_port, B1 => 
                           n455, B2 => REGISTERS_29_11_port, C1 => n466, C2 => 
                           REGISTERS_33_11_port, ZN => n14705);
   U13216 : OAI221_X1 port map( B1 => n11394, B2 => n477, C1 => n11522, C2 => 
                           n488, A => n14706, ZN => n14701);
   U13217 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_20_11_port, B1 => 
                           n510, B2 => REGISTERS_24_11_port, C1 => n521, C2 => 
                           REGISTERS_28_11_port, ZN => n14706);
   U13218 : OAI221_X1 port map( B1 => n11234, B2 => n532, C1 => n11362, C2 => 
                           n543, A => n14707, ZN => n14700);
   U13219 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_23_11_port, B1 => 
                           n565, B2 => REGISTERS_21_11_port, C1 => n576, C2 => 
                           REGISTERS_19_11_port, ZN => n14707);
   U13220 : NOR4_X1 port map( A1 => n14710, A2 => n14711, A3 => n14712, A4 => 
                           n14713, ZN => n14709);
   U13221 : OAI221_X1 port map( B1 => n11138, B2 => n312, C1 => n11074, C2 => 
                           n323, A => n14714, ZN => n14713);
   U13222 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_16_11_port, B1 => 
                           n119, B2 => REGISTERS_14_11_port, C1 => n13807, C2 
                           => REGISTERS_12_11_port, ZN => n14714);
   U13223 : OAI221_X1 port map( B1 => n11106, B2 => n13863, C1 => n10850, C2 =>
                           n13809, A => n14715, ZN => n14712);
   U13224 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_11_port, B1 => 
                           n13865, B2 => REGISTERS_9_11_port, C1 => n13813, C2 
                           => REGISTERS_7_11_port, ZN => n14715);
   U13225 : OAI221_X1 port map( B1 => n10946, B2 => n13866, C1 => n10690, C2 =>
                           n13815, A => n14716, ZN => n14711);
   U13226 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_11_port, B1 => 
                           n13868, B2 => REGISTERS_36_11_port, C1 => n13819, C2
                           => REGISTERS_3_11_port, ZN => n14716);
   U13227 : OAI221_X1 port map( B1 => n10786, B2 => n13869, C1 => n10658, C2 =>
                           n13821, A => n14717, ZN => n14710);
   U13228 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_11_port, B1 => 
                           n13871, B2 => REGISTERS_0_11_port, C1 => n13825, C2 
                           => REGISTERS_1_11_port, ZN => n14717);
   U13229 : NOR4_X1 port map( A1 => n14718, A2 => n14719, A3 => n14720, A4 => 
                           n14721, ZN => n14708);
   U13230 : OAI221_X1 port map( B1 => n11746, B2 => n367, C1 => n11010, C2 => 
                           n378, A => n14722, ZN => n14721);
   U13231 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_31_11_port, B1 => 
                           n400, B2 => REGISTERS_35_11_port, C1 => n411, C2 => 
                           REGISTERS_39_11_port, ZN => n14722);
   U13232 : OAI221_X1 port map( B1 => n11586, B2 => n422, C1 => n11714, C2 => 
                           n433, A => n14723, ZN => n14720);
   U13233 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_26_11_port, B1 => 
                           n455, B2 => REGISTERS_30_11_port, C1 => n466, C2 => 
                           REGISTERS_34_11_port, ZN => n14723);
   U13234 : OAI221_X1 port map( B1 => n11426, B2 => n477, C1 => n11554, C2 => 
                           n488, A => n14724, ZN => n14719);
   U13235 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_21_11_port, B1 => 
                           n510, B2 => REGISTERS_25_11_port, C1 => n521, C2 => 
                           REGISTERS_29_11_port, ZN => n14724);
   U13236 : OAI221_X1 port map( B1 => n11266, B2 => n532, C1 => n11394, C2 => 
                           n543, A => n14725, ZN => n14718);
   U13237 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_24_11_port, B1 => 
                           n565, B2 => REGISTERS_22_11_port, C1 => n576, C2 => 
                           REGISTERS_20_11_port, ZN => n14725);
   U13238 : AOI22_X1 port map( A1 => n13880, A2 => n4984, B1 => n13881, B2 => 
                           n4985, ZN => n14686);
   U13239 : NOR4_X1 port map( A1 => n14728, A2 => n14729, A3 => n14730, A4 => 
                           n14731, ZN => n14727);
   U13240 : OAI221_X1 port map( B1 => n11074, B2 => n312, C1 => n11010, C2 => 
                           n323, A => n14732, ZN => n14731);
   U13241 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_14_11_port, B1 => 
                           n13808, B2 => REGISTERS_38_11_port, C1 => n13889, C2
                           => REGISTERS_39_11_port, ZN => n14732);
   U13242 : OAI221_X1 port map( B1 => n10914, B2 => n13810, C1 => n10850, C2 =>
                           n13890, A => n14733, ZN => n14730);
   U13243 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_11_port, B1 => 
                           n343, B2 => REGISTERS_9_11_port, C1 => n13812, C2 =>
                           REGISTERS_16_11_port, ZN => n14733);
   U13244 : OAI221_X1 port map( B1 => n10754, B2 => n303, C1 => n10690, C2 => 
                           n13893, A => n14734, ZN => n14729);
   U13245 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_11_port, B1 => 
                           n354, B2 => REGISTERS_4_11_port, C1 => n13818, C2 =>
                           REGISTERS_11_11_port, ZN => n14734);
   U13246 : OAI221_X1 port map( B1 => n11618, B2 => n304, C1 => n10562, C2 => 
                           n13896, A => n14735, ZN => n14728);
   U13247 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_11_port, B1 => 
                           n13826, B2 => REGISTERS_0_11_port, C1 => n13824, C2 
                           => REGISTERS_6_11_port, ZN => n14735);
   U13248 : NOR4_X1 port map( A1 => n14736, A2 => n14737, A3 => n14738, A4 => 
                           n14739, ZN => n14726);
   U13249 : OAI221_X1 port map( B1 => n11682, B2 => n367, C1 => n10946, C2 => 
                           n378, A => n14740, ZN => n14739);
   U13250 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_29_11_port, B1 => 
                           n400, B2 => REGISTERS_33_11_port, C1 => n411, C2 => 
                           REGISTERS_37_11_port, ZN => n14740);
   U13251 : OAI221_X1 port map( B1 => n11522, B2 => n422, C1 => n11650, C2 => 
                           n433, A => n14741, ZN => n14738);
   U13252 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_24_11_port, B1 => 
                           n455, B2 => REGISTERS_28_11_port, C1 => n466, C2 => 
                           REGISTERS_32_11_port, ZN => n14741);
   U13253 : OAI221_X1 port map( B1 => n11362, B2 => n477, C1 => n11490, C2 => 
                           n488, A => n14742, ZN => n14737);
   U13254 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_19_11_port, B1 => 
                           n510, B2 => REGISTERS_23_11_port, C1 => n521, C2 => 
                           REGISTERS_27_11_port, ZN => n14742);
   U13255 : OAI221_X1 port map( B1 => n11202, B2 => n532, C1 => n11330, C2 => 
                           n543, A => n14743, ZN => n14736);
   U13256 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_22_11_port, B1 => 
                           n565, B2 => REGISTERS_20_11_port, C1 => n576, C2 => 
                           REGISTERS_18_11_port, ZN => n14743);
   U13257 : NOR4_X1 port map( A1 => n14746, A2 => n14747, A3 => n14748, A4 => 
                           n14749, ZN => n14745);
   U13258 : OAI221_X1 port map( B1 => n11042, B2 => n312, C1 => n10978, C2 => 
                           n323, A => n14750, ZN => n14749);
   U13259 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_13_11_port, B1 => 
                           n13808, B2 => REGISTERS_37_11_port, C1 => n13889, C2
                           => REGISTERS_38_11_port, ZN => n14750);
   U13260 : OAI221_X1 port map( B1 => n10882, B2 => n13810, C1 => n10818, C2 =>
                           n13890, A => n14751, ZN => n14748);
   U13261 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_11_port, B1 => 
                           n342, B2 => REGISTERS_8_11_port, C1 => n13812, C2 =>
                           REGISTERS_15_11_port, ZN => n14751);
   U13262 : OAI221_X1 port map( B1 => n10722, B2 => n303, C1 => n10658, C2 => 
                           n13893, A => n14752, ZN => n14747);
   U13263 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_11_port, B1 => 
                           n353, B2 => REGISTERS_3_11_port, C1 => n13818, C2 =>
                           REGISTERS_10_11_port, ZN => n14752);
   U13264 : OAI221_X1 port map( B1 => n11586, B2 => n304, C1 => n10508, C2 => 
                           n13896, A => n14753, ZN => n14746);
   U13265 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_11_port, B1 => 
                           n13917, B2 => REGISTERS_39_11_port, C1 => n13824, C2
                           => REGISTERS_5_11_port, ZN => n14753);
   U13266 : NOR4_X1 port map( A1 => n14754, A2 => n14755, A3 => n14756, A4 => 
                           n14757, ZN => n14744);
   U13267 : OAI221_X1 port map( B1 => n11650, B2 => n367, C1 => n10914, C2 => 
                           n378, A => n14758, ZN => n14757);
   U13268 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_28_11_port, B1 => 
                           n400, B2 => REGISTERS_32_11_port, C1 => n411, C2 => 
                           REGISTERS_36_11_port, ZN => n14758);
   U13269 : OAI221_X1 port map( B1 => n11490, B2 => n422, C1 => n11618, C2 => 
                           n433, A => n14759, ZN => n14756);
   U13270 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_23_11_port, B1 => 
                           n455, B2 => REGISTERS_27_11_port, C1 => n466, C2 => 
                           REGISTERS_31_11_port, ZN => n14759);
   U13271 : OAI221_X1 port map( B1 => n11330, B2 => n477, C1 => n11458, C2 => 
                           n488, A => n14760, ZN => n14755);
   U13272 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_18_11_port, B1 => 
                           n510, B2 => REGISTERS_22_11_port, C1 => n521, C2 => 
                           REGISTERS_26_11_port, ZN => n14760);
   U13273 : OAI221_X1 port map( B1 => n11170, B2 => n532, C1 => n11298, C2 => 
                           n543, A => n14761, ZN => n14754);
   U13274 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_21_11_port, B1 => 
                           n565, B2 => REGISTERS_19_11_port, C1 => n576, C2 => 
                           REGISTERS_17_11_port, ZN => n14761);
   U13275 : NAND3_X1 port map( A1 => n14762, A2 => n14763, A3 => n14764, ZN => 
                           n11892);
   U13276 : AOI221_X1 port map( B1 => n13792, B2 => n4989, C1 => n13793, C2 => 
                           MEM_IN(12), A => n14765, ZN => n14764);
   U13277 : OAI22_X1 port map( A1 => n10505, A2 => n251, B1 => n4991, B2 => 
                           n121, ZN => n14765);
   U13278 : NOR2_X1 port map( A1 => n5620, A2 => n13796, ZN => n5618);
   U13279 : INV_X1 port map( A => MEM_IN(12), ZN => n5620);
   U13280 : AOI22_X1 port map( A1 => n197, A2 => n4992, B1 => n150, B2 => n4993
                           , ZN => n14763);
   U13281 : NOR4_X1 port map( A1 => n14768, A2 => n14769, A3 => n14770, A4 => 
                           n14771, ZN => n14767);
   U13282 : OAI221_X1 port map( B1 => n11105, B2 => n312, C1 => n11041, C2 => 
                           n323, A => n14772, ZN => n14771);
   U13283 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_15_12_port, B1 => 
                           n13807, B2 => REGISTERS_11_12_port, C1 => n13808, C2
                           => REGISTERS_39_12_port, ZN => n14772);
   U13284 : OAI221_X1 port map( B1 => n10817, B2 => n13809, C1 => n10945, C2 =>
                           n13810, A => n14773, ZN => n14770);
   U13285 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_12_port, B1 =>
                           n13813, B2 => REGISTERS_6_12_port, C1 => n348, C2 =>
                           REGISTERS_10_12_port, ZN => n14773);
   U13286 : OAI221_X1 port map( B1 => n10657, B2 => n13815, C1 => n10785, C2 =>
                           n303, A => n14774, ZN => n14769);
   U13287 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_12_port, B1 =>
                           n13819, B2 => REGISTERS_2_12_port, C1 => n359, C2 =>
                           REGISTERS_5_12_port, ZN => n14774);
   U13288 : OAI221_X1 port map( B1 => n10625, B2 => n13821, C1 => n11649, C2 =>
                           n304, A => n14775, ZN => n14768);
   U13289 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_12_port, B1 => 
                           n13825, B2 => REGISTERS_0_12_port, C1 => n13826, C2 
                           => REGISTERS_1_12_port, ZN => n14775);
   U13290 : NOR4_X1 port map( A1 => n14776, A2 => n14777, A3 => n14778, A4 => 
                           n14779, ZN => n14766);
   U13291 : OAI221_X1 port map( B1 => n11713, B2 => n367, C1 => n10977, C2 => 
                           n378, A => n14780, ZN => n14779);
   U13292 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_30_12_port, B1 => 
                           n400, B2 => REGISTERS_34_12_port, C1 => n411, C2 => 
                           REGISTERS_38_12_port, ZN => n14780);
   U13293 : OAI221_X1 port map( B1 => n11553, B2 => n422, C1 => n11681, C2 => 
                           n433, A => n14781, ZN => n14778);
   U13294 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_25_12_port, B1 => 
                           n455, B2 => REGISTERS_29_12_port, C1 => n466, C2 => 
                           REGISTERS_33_12_port, ZN => n14781);
   U13295 : OAI221_X1 port map( B1 => n11393, B2 => n477, C1 => n11521, C2 => 
                           n488, A => n14782, ZN => n14777);
   U13296 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_20_12_port, B1 => 
                           n510, B2 => REGISTERS_24_12_port, C1 => n521, C2 => 
                           REGISTERS_28_12_port, ZN => n14782);
   U13297 : OAI221_X1 port map( B1 => n11233, B2 => n532, C1 => n11361, C2 => 
                           n543, A => n14783, ZN => n14776);
   U13298 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_23_12_port, B1 => 
                           n565, B2 => REGISTERS_21_12_port, C1 => n576, C2 => 
                           REGISTERS_19_12_port, ZN => n14783);
   U13299 : NOR4_X1 port map( A1 => n14786, A2 => n14787, A3 => n14788, A4 => 
                           n14789, ZN => n14785);
   U13300 : OAI221_X1 port map( B1 => n11137, B2 => n312, C1 => n11073, C2 => 
                           n323, A => n14790, ZN => n14789);
   U13301 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_16_12_port, B1 => 
                           n119, B2 => REGISTERS_14_12_port, C1 => n13807, C2 
                           => REGISTERS_12_12_port, ZN => n14790);
   U13302 : OAI221_X1 port map( B1 => n11105, B2 => n13863, C1 => n10849, C2 =>
                           n13809, A => n14791, ZN => n14788);
   U13303 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_12_port, B1 => 
                           n13865, B2 => REGISTERS_9_12_port, C1 => n13813, C2 
                           => REGISTERS_7_12_port, ZN => n14791);
   U13304 : OAI221_X1 port map( B1 => n10945, B2 => n13866, C1 => n10689, C2 =>
                           n13815, A => n14792, ZN => n14787);
   U13305 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_12_port, B1 => 
                           n13868, B2 => REGISTERS_36_12_port, C1 => n13819, C2
                           => REGISTERS_3_12_port, ZN => n14792);
   U13306 : OAI221_X1 port map( B1 => n10785, B2 => n13869, C1 => n10657, C2 =>
                           n13821, A => n14793, ZN => n14786);
   U13307 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_12_port, B1 => 
                           n13871, B2 => REGISTERS_0_12_port, C1 => n13825, C2 
                           => REGISTERS_1_12_port, ZN => n14793);
   U13308 : NOR4_X1 port map( A1 => n14794, A2 => n14795, A3 => n14796, A4 => 
                           n14797, ZN => n14784);
   U13309 : OAI221_X1 port map( B1 => n11745, B2 => n367, C1 => n11009, C2 => 
                           n378, A => n14798, ZN => n14797);
   U13310 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_31_12_port, B1 => 
                           n400, B2 => REGISTERS_35_12_port, C1 => n411, C2 => 
                           REGISTERS_39_12_port, ZN => n14798);
   U13311 : OAI221_X1 port map( B1 => n11585, B2 => n422, C1 => n11713, C2 => 
                           n433, A => n14799, ZN => n14796);
   U13312 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_26_12_port, B1 => 
                           n455, B2 => REGISTERS_30_12_port, C1 => n466, C2 => 
                           REGISTERS_34_12_port, ZN => n14799);
   U13313 : OAI221_X1 port map( B1 => n11425, B2 => n477, C1 => n11553, C2 => 
                           n488, A => n14800, ZN => n14795);
   U13314 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_21_12_port, B1 => 
                           n510, B2 => REGISTERS_25_12_port, C1 => n521, C2 => 
                           REGISTERS_29_12_port, ZN => n14800);
   U13315 : OAI221_X1 port map( B1 => n11265, B2 => n532, C1 => n11393, C2 => 
                           n543, A => n14801, ZN => n14794);
   U13316 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_24_12_port, B1 => 
                           n565, B2 => REGISTERS_22_12_port, C1 => n576, C2 => 
                           REGISTERS_20_12_port, ZN => n14801);
   U13317 : AOI22_X1 port map( A1 => n13880, A2 => n4994, B1 => n13881, B2 => 
                           n4995, ZN => n14762);
   U13318 : NOR4_X1 port map( A1 => n14804, A2 => n14805, A3 => n14806, A4 => 
                           n14807, ZN => n14803);
   U13319 : OAI221_X1 port map( B1 => n11073, B2 => n312, C1 => n11009, C2 => 
                           n323, A => n14808, ZN => n14807);
   U13320 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_14_12_port, B1 => 
                           n13808, B2 => REGISTERS_38_12_port, C1 => n13889, C2
                           => REGISTERS_39_12_port, ZN => n14808);
   U13321 : OAI221_X1 port map( B1 => n10913, B2 => n13810, C1 => n10849, C2 =>
                           n13890, A => n14809, ZN => n14806);
   U13322 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_12_port, B1 => 
                           n342, B2 => REGISTERS_9_12_port, C1 => n13812, C2 =>
                           REGISTERS_16_12_port, ZN => n14809);
   U13323 : OAI221_X1 port map( B1 => n10753, B2 => n303, C1 => n10689, C2 => 
                           n13893, A => n14810, ZN => n14805);
   U13324 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_12_port, B1 => 
                           n353, B2 => REGISTERS_4_12_port, C1 => n13818, C2 =>
                           REGISTERS_11_12_port, ZN => n14810);
   U13325 : OAI221_X1 port map( B1 => n11617, B2 => n304, C1 => n10561, C2 => 
                           n13896, A => n14811, ZN => n14804);
   U13326 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_12_port, B1 => 
                           n13826, B2 => REGISTERS_0_12_port, C1 => n13824, C2 
                           => REGISTERS_6_12_port, ZN => n14811);
   U13327 : NOR4_X1 port map( A1 => n14812, A2 => n14813, A3 => n14814, A4 => 
                           n14815, ZN => n14802);
   U13328 : OAI221_X1 port map( B1 => n11681, B2 => n367, C1 => n10945, C2 => 
                           n378, A => n14816, ZN => n14815);
   U13329 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_29_12_port, B1 => 
                           n400, B2 => REGISTERS_33_12_port, C1 => n411, C2 => 
                           REGISTERS_37_12_port, ZN => n14816);
   U13330 : OAI221_X1 port map( B1 => n11521, B2 => n422, C1 => n11649, C2 => 
                           n433, A => n14817, ZN => n14814);
   U13331 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_24_12_port, B1 => 
                           n455, B2 => REGISTERS_28_12_port, C1 => n466, C2 => 
                           REGISTERS_32_12_port, ZN => n14817);
   U13332 : OAI221_X1 port map( B1 => n11361, B2 => n477, C1 => n11489, C2 => 
                           n488, A => n14818, ZN => n14813);
   U13333 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_19_12_port, B1 => 
                           n510, B2 => REGISTERS_23_12_port, C1 => n521, C2 => 
                           REGISTERS_27_12_port, ZN => n14818);
   U13334 : OAI221_X1 port map( B1 => n11201, B2 => n532, C1 => n11329, C2 => 
                           n543, A => n14819, ZN => n14812);
   U13335 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_22_12_port, B1 => 
                           n565, B2 => REGISTERS_20_12_port, C1 => n576, C2 => 
                           REGISTERS_18_12_port, ZN => n14819);
   U13336 : NOR4_X1 port map( A1 => n14822, A2 => n14823, A3 => n14824, A4 => 
                           n14825, ZN => n14821);
   U13337 : OAI221_X1 port map( B1 => n11041, B2 => n312, C1 => n10977, C2 => 
                           n323, A => n14826, ZN => n14825);
   U13338 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_13_12_port, B1 => 
                           n13808, B2 => REGISTERS_37_12_port, C1 => n13889, C2
                           => REGISTERS_38_12_port, ZN => n14826);
   U13339 : OAI221_X1 port map( B1 => n10881, B2 => n13810, C1 => n10817, C2 =>
                           n13890, A => n14827, ZN => n14824);
   U13340 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_12_port, B1 => 
                           n342, B2 => REGISTERS_8_12_port, C1 => n13812, C2 =>
                           REGISTERS_15_12_port, ZN => n14827);
   U13341 : OAI221_X1 port map( B1 => n10721, B2 => n303, C1 => n10657, C2 => 
                           n13893, A => n14828, ZN => n14823);
   U13342 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_12_port, B1 => 
                           n353, B2 => REGISTERS_3_12_port, C1 => n13818, C2 =>
                           REGISTERS_10_12_port, ZN => n14828);
   U13343 : OAI221_X1 port map( B1 => n11585, B2 => n304, C1 => n10505, C2 => 
                           n13896, A => n14829, ZN => n14822);
   U13344 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_12_port, B1 => 
                           n13917, B2 => REGISTERS_39_12_port, C1 => n13824, C2
                           => REGISTERS_5_12_port, ZN => n14829);
   U13345 : NOR4_X1 port map( A1 => n14830, A2 => n14831, A3 => n14832, A4 => 
                           n14833, ZN => n14820);
   U13346 : OAI221_X1 port map( B1 => n11649, B2 => n367, C1 => n10913, C2 => 
                           n378, A => n14834, ZN => n14833);
   U13347 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_28_12_port, B1 => 
                           n400, B2 => REGISTERS_32_12_port, C1 => n411, C2 => 
                           REGISTERS_36_12_port, ZN => n14834);
   U13348 : OAI221_X1 port map( B1 => n11489, B2 => n422, C1 => n11617, C2 => 
                           n433, A => n14835, ZN => n14832);
   U13349 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_23_12_port, B1 => 
                           n455, B2 => REGISTERS_27_12_port, C1 => n466, C2 => 
                           REGISTERS_31_12_port, ZN => n14835);
   U13350 : OAI221_X1 port map( B1 => n11329, B2 => n477, C1 => n11457, C2 => 
                           n488, A => n14836, ZN => n14831);
   U13351 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_18_12_port, B1 => 
                           n510, B2 => REGISTERS_22_12_port, C1 => n521, C2 => 
                           REGISTERS_26_12_port, ZN => n14836);
   U13352 : OAI221_X1 port map( B1 => n11169, B2 => n532, C1 => n11297, C2 => 
                           n543, A => n14837, ZN => n14830);
   U13353 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_21_12_port, B1 => 
                           n565, B2 => REGISTERS_19_12_port, C1 => n576, C2 => 
                           REGISTERS_17_12_port, ZN => n14837);
   U13354 : NAND3_X1 port map( A1 => n14838, A2 => n14839, A3 => n14840, ZN => 
                           n11891);
   U13355 : AOI221_X1 port map( B1 => n13792, B2 => n4999, C1 => n13793, C2 => 
                           MEM_IN(13), A => n14841, ZN => n14840);
   U13356 : OAI22_X1 port map( A1 => n10502, A2 => n251, B1 => n5001, B2 => 
                           n121, ZN => n14841);
   U13357 : NOR2_X1 port map( A1 => n5627, A2 => n13796, ZN => n5625);
   U13358 : INV_X1 port map( A => MEM_IN(13), ZN => n5627);
   U13359 : AOI22_X1 port map( A1 => n197, A2 => n5002, B1 => n150, B2 => n5003
                           , ZN => n14839);
   U13360 : NOR4_X1 port map( A1 => n14844, A2 => n14845, A3 => n14846, A4 => 
                           n14847, ZN => n14843);
   U13361 : OAI221_X1 port map( B1 => n11104, B2 => n312, C1 => n11040, C2 => 
                           n323, A => n14848, ZN => n14847);
   U13362 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_15_13_port, B1 => 
                           n13807, B2 => REGISTERS_11_13_port, C1 => n13808, C2
                           => REGISTERS_39_13_port, ZN => n14848);
   U13363 : OAI221_X1 port map( B1 => n10816, B2 => n13809, C1 => n10944, C2 =>
                           n13810, A => n14849, ZN => n14846);
   U13364 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_13_port, B1 =>
                           n13813, B2 => REGISTERS_6_13_port, C1 => n348, C2 =>
                           REGISTERS_10_13_port, ZN => n14849);
   U13365 : OAI221_X1 port map( B1 => n10656, B2 => n13815, C1 => n10784, C2 =>
                           n303, A => n14850, ZN => n14845);
   U13366 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_13_port, B1 =>
                           n13819, B2 => REGISTERS_2_13_port, C1 => n359, C2 =>
                           REGISTERS_5_13_port, ZN => n14850);
   U13367 : OAI221_X1 port map( B1 => n10624, B2 => n13821, C1 => n11648, C2 =>
                           n304, A => n14851, ZN => n14844);
   U13368 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_13_port, B1 => 
                           n13825, B2 => REGISTERS_0_13_port, C1 => n13826, C2 
                           => REGISTERS_1_13_port, ZN => n14851);
   U13369 : NOR4_X1 port map( A1 => n14852, A2 => n14853, A3 => n14854, A4 => 
                           n14855, ZN => n14842);
   U13370 : OAI221_X1 port map( B1 => n11712, B2 => n367, C1 => n10976, C2 => 
                           n378, A => n14856, ZN => n14855);
   U13371 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_30_13_port, B1 => 
                           n400, B2 => REGISTERS_34_13_port, C1 => n411, C2 => 
                           REGISTERS_38_13_port, ZN => n14856);
   U13372 : OAI221_X1 port map( B1 => n11552, B2 => n422, C1 => n11680, C2 => 
                           n433, A => n14857, ZN => n14854);
   U13373 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_25_13_port, B1 => 
                           n455, B2 => REGISTERS_29_13_port, C1 => n466, C2 => 
                           REGISTERS_33_13_port, ZN => n14857);
   U13374 : OAI221_X1 port map( B1 => n11392, B2 => n477, C1 => n11520, C2 => 
                           n488, A => n14858, ZN => n14853);
   U13375 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_20_13_port, B1 => 
                           n510, B2 => REGISTERS_24_13_port, C1 => n521, C2 => 
                           REGISTERS_28_13_port, ZN => n14858);
   U13376 : OAI221_X1 port map( B1 => n11232, B2 => n532, C1 => n11360, C2 => 
                           n543, A => n14859, ZN => n14852);
   U13377 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_23_13_port, B1 => 
                           n565, B2 => REGISTERS_21_13_port, C1 => n576, C2 => 
                           REGISTERS_19_13_port, ZN => n14859);
   U13378 : NOR4_X1 port map( A1 => n14862, A2 => n14863, A3 => n14864, A4 => 
                           n14865, ZN => n14861);
   U13379 : OAI221_X1 port map( B1 => n11136, B2 => n312, C1 => n11072, C2 => 
                           n323, A => n14866, ZN => n14865);
   U13380 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_16_13_port, B1 => 
                           n119, B2 => REGISTERS_14_13_port, C1 => n13807, C2 
                           => REGISTERS_12_13_port, ZN => n14866);
   U13381 : OAI221_X1 port map( B1 => n11104, B2 => n13863, C1 => n10848, C2 =>
                           n13809, A => n14867, ZN => n14864);
   U13382 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_13_port, B1 => 
                           n13865, B2 => REGISTERS_9_13_port, C1 => n13813, C2 
                           => REGISTERS_7_13_port, ZN => n14867);
   U13383 : OAI221_X1 port map( B1 => n10944, B2 => n13866, C1 => n10688, C2 =>
                           n13815, A => n14868, ZN => n14863);
   U13384 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_13_port, B1 => 
                           n13868, B2 => REGISTERS_36_13_port, C1 => n13819, C2
                           => REGISTERS_3_13_port, ZN => n14868);
   U13385 : OAI221_X1 port map( B1 => n10784, B2 => n13869, C1 => n10656, C2 =>
                           n13821, A => n14869, ZN => n14862);
   U13386 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_13_port, B1 => 
                           n13871, B2 => REGISTERS_0_13_port, C1 => n13825, C2 
                           => REGISTERS_1_13_port, ZN => n14869);
   U13387 : NOR4_X1 port map( A1 => n14870, A2 => n14871, A3 => n14872, A4 => 
                           n14873, ZN => n14860);
   U13388 : OAI221_X1 port map( B1 => n11744, B2 => n367, C1 => n11008, C2 => 
                           n378, A => n14874, ZN => n14873);
   U13389 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_31_13_port, B1 => 
                           n400, B2 => REGISTERS_35_13_port, C1 => n411, C2 => 
                           REGISTERS_39_13_port, ZN => n14874);
   U13390 : OAI221_X1 port map( B1 => n11584, B2 => n422, C1 => n11712, C2 => 
                           n433, A => n14875, ZN => n14872);
   U13391 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_26_13_port, B1 => 
                           n455, B2 => REGISTERS_30_13_port, C1 => n466, C2 => 
                           REGISTERS_34_13_port, ZN => n14875);
   U13392 : OAI221_X1 port map( B1 => n11424, B2 => n477, C1 => n11552, C2 => 
                           n488, A => n14876, ZN => n14871);
   U13393 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_21_13_port, B1 => 
                           n510, B2 => REGISTERS_25_13_port, C1 => n521, C2 => 
                           REGISTERS_29_13_port, ZN => n14876);
   U13394 : OAI221_X1 port map( B1 => n11264, B2 => n532, C1 => n11392, C2 => 
                           n543, A => n14877, ZN => n14870);
   U13395 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_24_13_port, B1 => 
                           n565, B2 => REGISTERS_22_13_port, C1 => n576, C2 => 
                           REGISTERS_20_13_port, ZN => n14877);
   U13396 : AOI22_X1 port map( A1 => n13880, A2 => n5004, B1 => n13881, B2 => 
                           n5005, ZN => n14838);
   U13397 : NOR4_X1 port map( A1 => n14880, A2 => n14881, A3 => n14882, A4 => 
                           n14883, ZN => n14879);
   U13398 : OAI221_X1 port map( B1 => n11072, B2 => n312, C1 => n11008, C2 => 
                           n323, A => n14884, ZN => n14883);
   U13399 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_14_13_port, B1 => 
                           n13808, B2 => REGISTERS_38_13_port, C1 => n13889, C2
                           => REGISTERS_39_13_port, ZN => n14884);
   U13400 : OAI221_X1 port map( B1 => n10912, B2 => n13810, C1 => n10848, C2 =>
                           n13890, A => n14885, ZN => n14882);
   U13401 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_13_port, B1 => 
                           n343, B2 => REGISTERS_9_13_port, C1 => n13812, C2 =>
                           REGISTERS_16_13_port, ZN => n14885);
   U13402 : OAI221_X1 port map( B1 => n10752, B2 => n303, C1 => n10688, C2 => 
                           n13893, A => n14886, ZN => n14881);
   U13403 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_13_port, B1 => 
                           n354, B2 => REGISTERS_4_13_port, C1 => n13818, C2 =>
                           REGISTERS_11_13_port, ZN => n14886);
   U13404 : OAI221_X1 port map( B1 => n11616, B2 => n304, C1 => n10560, C2 => 
                           n13896, A => n14887, ZN => n14880);
   U13405 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_13_port, B1 => 
                           n13826, B2 => REGISTERS_0_13_port, C1 => n13824, C2 
                           => REGISTERS_6_13_port, ZN => n14887);
   U13406 : NOR4_X1 port map( A1 => n14888, A2 => n14889, A3 => n14890, A4 => 
                           n14891, ZN => n14878);
   U13407 : OAI221_X1 port map( B1 => n11680, B2 => n367, C1 => n10944, C2 => 
                           n378, A => n14892, ZN => n14891);
   U13408 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_29_13_port, B1 => 
                           n400, B2 => REGISTERS_33_13_port, C1 => n411, C2 => 
                           REGISTERS_37_13_port, ZN => n14892);
   U13409 : OAI221_X1 port map( B1 => n11520, B2 => n422, C1 => n11648, C2 => 
                           n433, A => n14893, ZN => n14890);
   U13410 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_24_13_port, B1 => 
                           n455, B2 => REGISTERS_28_13_port, C1 => n466, C2 => 
                           REGISTERS_32_13_port, ZN => n14893);
   U13411 : OAI221_X1 port map( B1 => n11360, B2 => n477, C1 => n11488, C2 => 
                           n488, A => n14894, ZN => n14889);
   U13412 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_19_13_port, B1 => 
                           n510, B2 => REGISTERS_23_13_port, C1 => n521, C2 => 
                           REGISTERS_27_13_port, ZN => n14894);
   U13413 : OAI221_X1 port map( B1 => n11200, B2 => n532, C1 => n11328, C2 => 
                           n543, A => n14895, ZN => n14888);
   U13414 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_22_13_port, B1 => 
                           n565, B2 => REGISTERS_20_13_port, C1 => n576, C2 => 
                           REGISTERS_18_13_port, ZN => n14895);
   U13415 : NOR4_X1 port map( A1 => n14898, A2 => n14899, A3 => n14900, A4 => 
                           n14901, ZN => n14897);
   U13416 : OAI221_X1 port map( B1 => n11040, B2 => n312, C1 => n10976, C2 => 
                           n323, A => n14902, ZN => n14901);
   U13417 : AOI222_X1 port map( A1 => n334, A2 => REGISTERS_13_13_port, B1 => 
                           n13808, B2 => REGISTERS_37_13_port, C1 => n13889, C2
                           => REGISTERS_38_13_port, ZN => n14902);
   U13418 : OAI221_X1 port map( B1 => n10880, B2 => n13810, C1 => n10816, C2 =>
                           n13890, A => n14903, ZN => n14900);
   U13419 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_13_port, B1 => 
                           n343, B2 => REGISTERS_8_13_port, C1 => n13812, C2 =>
                           REGISTERS_15_13_port, ZN => n14903);
   U13420 : OAI221_X1 port map( B1 => n10720, B2 => n303, C1 => n10656, C2 => 
                           n13893, A => n14904, ZN => n14899);
   U13421 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_13_port, B1 => 
                           n354, B2 => REGISTERS_3_13_port, C1 => n13818, C2 =>
                           REGISTERS_10_13_port, ZN => n14904);
   U13422 : OAI221_X1 port map( B1 => n11584, B2 => n304, C1 => n10502, C2 => 
                           n13896, A => n14905, ZN => n14898);
   U13423 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_13_port, B1 => 
                           n13917, B2 => REGISTERS_39_13_port, C1 => n13824, C2
                           => REGISTERS_5_13_port, ZN => n14905);
   U13424 : NOR4_X1 port map( A1 => n14906, A2 => n14907, A3 => n14908, A4 => 
                           n14909, ZN => n14896);
   U13425 : OAI221_X1 port map( B1 => n11648, B2 => n367, C1 => n10912, C2 => 
                           n378, A => n14910, ZN => n14909);
   U13426 : AOI222_X1 port map( A1 => n389, A2 => REGISTERS_28_13_port, B1 => 
                           n400, B2 => REGISTERS_32_13_port, C1 => n411, C2 => 
                           REGISTERS_36_13_port, ZN => n14910);
   U13427 : OAI221_X1 port map( B1 => n11488, B2 => n422, C1 => n11616, C2 => 
                           n433, A => n14911, ZN => n14908);
   U13428 : AOI222_X1 port map( A1 => n444, A2 => REGISTERS_23_13_port, B1 => 
                           n455, B2 => REGISTERS_27_13_port, C1 => n466, C2 => 
                           REGISTERS_31_13_port, ZN => n14911);
   U13429 : OAI221_X1 port map( B1 => n11328, B2 => n477, C1 => n11456, C2 => 
                           n488, A => n14912, ZN => n14907);
   U13430 : AOI222_X1 port map( A1 => n499, A2 => REGISTERS_18_13_port, B1 => 
                           n510, B2 => REGISTERS_22_13_port, C1 => n521, C2 => 
                           REGISTERS_26_13_port, ZN => n14912);
   U13431 : OAI221_X1 port map( B1 => n11168, B2 => n532, C1 => n11296, C2 => 
                           n543, A => n14913, ZN => n14906);
   U13432 : AOI222_X1 port map( A1 => n554, A2 => REGISTERS_21_13_port, B1 => 
                           n565, B2 => REGISTERS_19_13_port, C1 => n576, C2 => 
                           REGISTERS_17_13_port, ZN => n14913);
   U13433 : NAND3_X1 port map( A1 => n14914, A2 => n14915, A3 => n14916, ZN => 
                           n11890);
   U13434 : AOI221_X1 port map( B1 => n13792, B2 => n5009, C1 => n13793, C2 => 
                           MEM_IN(14), A => n14917, ZN => n14916);
   U13435 : OAI22_X1 port map( A1 => n10499, A2 => n251, B1 => n5011, B2 => 
                           n121, ZN => n14917);
   U13436 : NOR2_X1 port map( A1 => n5634, A2 => n13796, ZN => n5632);
   U13437 : INV_X1 port map( A => MEM_IN(14), ZN => n5634);
   U13438 : AOI22_X1 port map( A1 => n197, A2 => n5012, B1 => n150, B2 => n5013
                           , ZN => n14915);
   U13439 : NOR4_X1 port map( A1 => n14920, A2 => n14921, A3 => n14922, A4 => 
                           n14923, ZN => n14919);
   U13440 : OAI221_X1 port map( B1 => n11103, B2 => n311, C1 => n11039, C2 => 
                           n322, A => n14924, ZN => n14923);
   U13441 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_15_14_port, B1 => 
                           n13807, B2 => REGISTERS_11_14_port, C1 => n13808, C2
                           => REGISTERS_39_14_port, ZN => n14924);
   U13442 : OAI221_X1 port map( B1 => n10815, B2 => n13809, C1 => n10943, C2 =>
                           n13810, A => n14925, ZN => n14922);
   U13443 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_14_port, B1 =>
                           n13813, B2 => REGISTERS_6_14_port, C1 => n348, C2 =>
                           REGISTERS_10_14_port, ZN => n14925);
   U13444 : OAI221_X1 port map( B1 => n10655, B2 => n13815, C1 => n10783, C2 =>
                           n303, A => n14926, ZN => n14921);
   U13445 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_14_port, B1 =>
                           n13819, B2 => REGISTERS_2_14_port, C1 => n359, C2 =>
                           REGISTERS_5_14_port, ZN => n14926);
   U13446 : OAI221_X1 port map( B1 => n10623, B2 => n13821, C1 => n11647, C2 =>
                           n304, A => n14927, ZN => n14920);
   U13447 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_14_port, B1 => 
                           n13825, B2 => REGISTERS_0_14_port, C1 => n13826, C2 
                           => REGISTERS_1_14_port, ZN => n14927);
   U13448 : NOR4_X1 port map( A1 => n14928, A2 => n14929, A3 => n14930, A4 => 
                           n14931, ZN => n14918);
   U13449 : OAI221_X1 port map( B1 => n11711, B2 => n366, C1 => n10975, C2 => 
                           n378, A => n14932, ZN => n14931);
   U13450 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_30_14_port, B1 => 
                           n399, B2 => REGISTERS_34_14_port, C1 => n410, C2 => 
                           REGISTERS_38_14_port, ZN => n14932);
   U13451 : OAI221_X1 port map( B1 => n11551, B2 => n421, C1 => n11679, C2 => 
                           n432, A => n14933, ZN => n14930);
   U13452 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_25_14_port, B1 => 
                           n454, B2 => REGISTERS_29_14_port, C1 => n465, C2 => 
                           REGISTERS_33_14_port, ZN => n14933);
   U13453 : OAI221_X1 port map( B1 => n11391, B2 => n476, C1 => n11519, C2 => 
                           n487, A => n14934, ZN => n14929);
   U13454 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_20_14_port, B1 => 
                           n509, B2 => REGISTERS_24_14_port, C1 => n520, C2 => 
                           REGISTERS_28_14_port, ZN => n14934);
   U13455 : OAI221_X1 port map( B1 => n11231, B2 => n531, C1 => n11359, C2 => 
                           n542, A => n14935, ZN => n14928);
   U13456 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_23_14_port, B1 => 
                           n564, B2 => REGISTERS_21_14_port, C1 => n575, C2 => 
                           REGISTERS_19_14_port, ZN => n14935);
   U13457 : NOR4_X1 port map( A1 => n14938, A2 => n14939, A3 => n14940, A4 => 
                           n14941, ZN => n14937);
   U13458 : OAI221_X1 port map( B1 => n11135, B2 => n311, C1 => n11071, C2 => 
                           n322, A => n14942, ZN => n14941);
   U13459 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_16_14_port, B1 => 
                           n119, B2 => REGISTERS_14_14_port, C1 => n13807, C2 
                           => REGISTERS_12_14_port, ZN => n14942);
   U13460 : OAI221_X1 port map( B1 => n11103, B2 => n13863, C1 => n10847, C2 =>
                           n13809, A => n14943, ZN => n14940);
   U13461 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_14_port, B1 => 
                           n13865, B2 => REGISTERS_9_14_port, C1 => n13813, C2 
                           => REGISTERS_7_14_port, ZN => n14943);
   U13462 : OAI221_X1 port map( B1 => n10943, B2 => n13866, C1 => n10687, C2 =>
                           n13815, A => n14944, ZN => n14939);
   U13463 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_14_port, B1 => 
                           n13868, B2 => REGISTERS_36_14_port, C1 => n13819, C2
                           => REGISTERS_3_14_port, ZN => n14944);
   U13464 : OAI221_X1 port map( B1 => n10783, B2 => n13869, C1 => n10655, C2 =>
                           n13821, A => n14945, ZN => n14938);
   U13465 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_14_port, B1 => 
                           n13871, B2 => REGISTERS_0_14_port, C1 => n13825, C2 
                           => REGISTERS_1_14_port, ZN => n14945);
   U13466 : NOR4_X1 port map( A1 => n14946, A2 => n14947, A3 => n14948, A4 => 
                           n14949, ZN => n14936);
   U13467 : OAI221_X1 port map( B1 => n11743, B2 => n366, C1 => n11007, C2 => 
                           n377, A => n14950, ZN => n14949);
   U13468 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_31_14_port, B1 => 
                           n399, B2 => REGISTERS_35_14_port, C1 => n410, C2 => 
                           REGISTERS_39_14_port, ZN => n14950);
   U13469 : OAI221_X1 port map( B1 => n11583, B2 => n421, C1 => n11711, C2 => 
                           n432, A => n14951, ZN => n14948);
   U13470 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_26_14_port, B1 => 
                           n454, B2 => REGISTERS_30_14_port, C1 => n465, C2 => 
                           REGISTERS_34_14_port, ZN => n14951);
   U13471 : OAI221_X1 port map( B1 => n11423, B2 => n476, C1 => n11551, C2 => 
                           n487, A => n14952, ZN => n14947);
   U13472 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_21_14_port, B1 => 
                           n509, B2 => REGISTERS_25_14_port, C1 => n520, C2 => 
                           REGISTERS_29_14_port, ZN => n14952);
   U13473 : OAI221_X1 port map( B1 => n11263, B2 => n531, C1 => n11391, C2 => 
                           n542, A => n14953, ZN => n14946);
   U13474 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_24_14_port, B1 => 
                           n564, B2 => REGISTERS_22_14_port, C1 => n575, C2 => 
                           REGISTERS_20_14_port, ZN => n14953);
   U13475 : AOI22_X1 port map( A1 => n13880, A2 => n5014, B1 => n13881, B2 => 
                           n5015, ZN => n14914);
   U13476 : NOR4_X1 port map( A1 => n14956, A2 => n14957, A3 => n14958, A4 => 
                           n14959, ZN => n14955);
   U13477 : OAI221_X1 port map( B1 => n11071, B2 => n311, C1 => n11007, C2 => 
                           n322, A => n14960, ZN => n14959);
   U13478 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_14_14_port, B1 => 
                           n13808, B2 => REGISTERS_38_14_port, C1 => n13889, C2
                           => REGISTERS_39_14_port, ZN => n14960);
   U13479 : OAI221_X1 port map( B1 => n10911, B2 => n13810, C1 => n10847, C2 =>
                           n13890, A => n14961, ZN => n14958);
   U13480 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_14_port, B1 => 
                           n343, B2 => REGISTERS_9_14_port, C1 => n13812, C2 =>
                           REGISTERS_16_14_port, ZN => n14961);
   U13481 : OAI221_X1 port map( B1 => n10751, B2 => n303, C1 => n10687, C2 => 
                           n13893, A => n14962, ZN => n14957);
   U13482 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_14_port, B1 => 
                           n354, B2 => REGISTERS_4_14_port, C1 => n13818, C2 =>
                           REGISTERS_11_14_port, ZN => n14962);
   U13483 : OAI221_X1 port map( B1 => n11615, B2 => n304, C1 => n10559, C2 => 
                           n13896, A => n14963, ZN => n14956);
   U13484 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_14_port, B1 => 
                           n13826, B2 => REGISTERS_0_14_port, C1 => n13824, C2 
                           => REGISTERS_6_14_port, ZN => n14963);
   U13485 : NOR4_X1 port map( A1 => n14964, A2 => n14965, A3 => n14966, A4 => 
                           n14967, ZN => n14954);
   U13486 : OAI221_X1 port map( B1 => n11679, B2 => n366, C1 => n10943, C2 => 
                           n377, A => n14968, ZN => n14967);
   U13487 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_29_14_port, B1 => 
                           n399, B2 => REGISTERS_33_14_port, C1 => n410, C2 => 
                           REGISTERS_37_14_port, ZN => n14968);
   U13488 : OAI221_X1 port map( B1 => n11519, B2 => n421, C1 => n11647, C2 => 
                           n432, A => n14969, ZN => n14966);
   U13489 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_24_14_port, B1 => 
                           n454, B2 => REGISTERS_28_14_port, C1 => n465, C2 => 
                           REGISTERS_32_14_port, ZN => n14969);
   U13490 : OAI221_X1 port map( B1 => n11359, B2 => n476, C1 => n11487, C2 => 
                           n487, A => n14970, ZN => n14965);
   U13491 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_19_14_port, B1 => 
                           n509, B2 => REGISTERS_23_14_port, C1 => n520, C2 => 
                           REGISTERS_27_14_port, ZN => n14970);
   U13492 : OAI221_X1 port map( B1 => n11199, B2 => n531, C1 => n11327, C2 => 
                           n542, A => n14971, ZN => n14964);
   U13493 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_22_14_port, B1 => 
                           n564, B2 => REGISTERS_20_14_port, C1 => n575, C2 => 
                           REGISTERS_18_14_port, ZN => n14971);
   U13494 : NOR4_X1 port map( A1 => n14974, A2 => n14975, A3 => n14976, A4 => 
                           n14977, ZN => n14973);
   U13495 : OAI221_X1 port map( B1 => n11039, B2 => n311, C1 => n10975, C2 => 
                           n322, A => n14978, ZN => n14977);
   U13496 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_13_14_port, B1 => 
                           n13808, B2 => REGISTERS_37_14_port, C1 => n13889, C2
                           => REGISTERS_38_14_port, ZN => n14978);
   U13497 : OAI221_X1 port map( B1 => n10879, B2 => n13810, C1 => n10815, C2 =>
                           n13890, A => n14979, ZN => n14976);
   U13498 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_14_port, B1 => 
                           n343, B2 => REGISTERS_8_14_port, C1 => n13812, C2 =>
                           REGISTERS_15_14_port, ZN => n14979);
   U13499 : OAI221_X1 port map( B1 => n10719, B2 => n303, C1 => n10655, C2 => 
                           n13893, A => n14980, ZN => n14975);
   U13500 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_14_port, B1 => 
                           n354, B2 => REGISTERS_3_14_port, C1 => n13818, C2 =>
                           REGISTERS_10_14_port, ZN => n14980);
   U13501 : OAI221_X1 port map( B1 => n11583, B2 => n304, C1 => n10499, C2 => 
                           n13896, A => n14981, ZN => n14974);
   U13502 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_14_port, B1 => 
                           n13917, B2 => REGISTERS_39_14_port, C1 => n13824, C2
                           => REGISTERS_5_14_port, ZN => n14981);
   U13503 : NOR4_X1 port map( A1 => n14982, A2 => n14983, A3 => n14984, A4 => 
                           n14985, ZN => n14972);
   U13504 : OAI221_X1 port map( B1 => n11647, B2 => n366, C1 => n10911, C2 => 
                           n377, A => n14986, ZN => n14985);
   U13505 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_28_14_port, B1 => 
                           n399, B2 => REGISTERS_32_14_port, C1 => n410, C2 => 
                           REGISTERS_36_14_port, ZN => n14986);
   U13506 : OAI221_X1 port map( B1 => n11487, B2 => n421, C1 => n11615, C2 => 
                           n432, A => n14987, ZN => n14984);
   U13507 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_23_14_port, B1 => 
                           n454, B2 => REGISTERS_27_14_port, C1 => n465, C2 => 
                           REGISTERS_31_14_port, ZN => n14987);
   U13508 : OAI221_X1 port map( B1 => n11327, B2 => n476, C1 => n11455, C2 => 
                           n487, A => n14988, ZN => n14983);
   U13509 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_18_14_port, B1 => 
                           n509, B2 => REGISTERS_22_14_port, C1 => n520, C2 => 
                           REGISTERS_26_14_port, ZN => n14988);
   U13510 : OAI221_X1 port map( B1 => n11167, B2 => n531, C1 => n11295, C2 => 
                           n542, A => n14989, ZN => n14982);
   U13511 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_21_14_port, B1 => 
                           n564, B2 => REGISTERS_19_14_port, C1 => n575, C2 => 
                           REGISTERS_17_14_port, ZN => n14989);
   U13512 : NAND3_X1 port map( A1 => n14990, A2 => n14991, A3 => n14992, ZN => 
                           n11889);
   U13513 : AOI221_X1 port map( B1 => n13792, B2 => n5019, C1 => n13793, C2 => 
                           MEM_IN(15), A => n14993, ZN => n14992);
   U13514 : OAI22_X1 port map( A1 => n10496, A2 => n251, B1 => n5021, B2 => 
                           n121, ZN => n14993);
   U13515 : NOR2_X1 port map( A1 => n5641, A2 => n13796, ZN => n5639);
   U13516 : INV_X1 port map( A => MEM_IN(15), ZN => n5641);
   U13517 : AOI22_X1 port map( A1 => n197, A2 => n5022, B1 => n150, B2 => n5023
                           , ZN => n14991);
   U13518 : NOR4_X1 port map( A1 => n14996, A2 => n14997, A3 => n14998, A4 => 
                           n14999, ZN => n14995);
   U13519 : OAI221_X1 port map( B1 => n11102, B2 => n311, C1 => n11038, C2 => 
                           n322, A => n15000, ZN => n14999);
   U13520 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_15_15_port, B1 => 
                           n13807, B2 => REGISTERS_11_15_port, C1 => n13808, C2
                           => REGISTERS_39_15_port, ZN => n15000);
   U13521 : OAI221_X1 port map( B1 => n10814, B2 => n13809, C1 => n10942, C2 =>
                           n13810, A => n15001, ZN => n14998);
   U13522 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_15_port, B1 =>
                           n13813, B2 => REGISTERS_6_15_port, C1 => n348, C2 =>
                           REGISTERS_10_15_port, ZN => n15001);
   U13523 : OAI221_X1 port map( B1 => n10654, B2 => n13815, C1 => n10782, C2 =>
                           n303, A => n15002, ZN => n14997);
   U13524 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_15_port, B1 =>
                           n13819, B2 => REGISTERS_2_15_port, C1 => n359, C2 =>
                           REGISTERS_5_15_port, ZN => n15002);
   U13525 : OAI221_X1 port map( B1 => n10622, B2 => n13821, C1 => n11646, C2 =>
                           n304, A => n15003, ZN => n14996);
   U13526 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_15_port, B1 => 
                           n13825, B2 => REGISTERS_0_15_port, C1 => n13826, C2 
                           => REGISTERS_1_15_port, ZN => n15003);
   U13527 : NOR4_X1 port map( A1 => n15004, A2 => n15005, A3 => n15006, A4 => 
                           n15007, ZN => n14994);
   U13528 : OAI221_X1 port map( B1 => n11710, B2 => n366, C1 => n10974, C2 => 
                           n377, A => n15008, ZN => n15007);
   U13529 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_30_15_port, B1 => 
                           n399, B2 => REGISTERS_34_15_port, C1 => n410, C2 => 
                           REGISTERS_38_15_port, ZN => n15008);
   U13530 : OAI221_X1 port map( B1 => n11550, B2 => n421, C1 => n11678, C2 => 
                           n432, A => n15009, ZN => n15006);
   U13531 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_25_15_port, B1 => 
                           n454, B2 => REGISTERS_29_15_port, C1 => n465, C2 => 
                           REGISTERS_33_15_port, ZN => n15009);
   U13532 : OAI221_X1 port map( B1 => n11390, B2 => n476, C1 => n11518, C2 => 
                           n487, A => n15010, ZN => n15005);
   U13533 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_20_15_port, B1 => 
                           n509, B2 => REGISTERS_24_15_port, C1 => n520, C2 => 
                           REGISTERS_28_15_port, ZN => n15010);
   U13534 : OAI221_X1 port map( B1 => n11230, B2 => n531, C1 => n11358, C2 => 
                           n542, A => n15011, ZN => n15004);
   U13535 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_23_15_port, B1 => 
                           n564, B2 => REGISTERS_21_15_port, C1 => n575, C2 => 
                           REGISTERS_19_15_port, ZN => n15011);
   U13536 : NOR4_X1 port map( A1 => n15014, A2 => n15015, A3 => n15016, A4 => 
                           n15017, ZN => n15013);
   U13537 : OAI221_X1 port map( B1 => n11134, B2 => n311, C1 => n11070, C2 => 
                           n322, A => n15018, ZN => n15017);
   U13538 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_16_15_port, B1 => 
                           n119, B2 => REGISTERS_14_15_port, C1 => n13807, C2 
                           => REGISTERS_12_15_port, ZN => n15018);
   U13539 : OAI221_X1 port map( B1 => n11102, B2 => n13863, C1 => n10846, C2 =>
                           n13809, A => n15019, ZN => n15016);
   U13540 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_15_port, B1 => 
                           n13865, B2 => REGISTERS_9_15_port, C1 => n13813, C2 
                           => REGISTERS_7_15_port, ZN => n15019);
   U13541 : OAI221_X1 port map( B1 => n10942, B2 => n13866, C1 => n10686, C2 =>
                           n13815, A => n15020, ZN => n15015);
   U13542 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_15_port, B1 => 
                           n13868, B2 => REGISTERS_36_15_port, C1 => n13819, C2
                           => REGISTERS_3_15_port, ZN => n15020);
   U13543 : OAI221_X1 port map( B1 => n10782, B2 => n13869, C1 => n10654, C2 =>
                           n13821, A => n15021, ZN => n15014);
   U13544 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_15_port, B1 => 
                           n13871, B2 => REGISTERS_0_15_port, C1 => n13825, C2 
                           => REGISTERS_1_15_port, ZN => n15021);
   U13545 : NOR4_X1 port map( A1 => n15022, A2 => n15023, A3 => n15024, A4 => 
                           n15025, ZN => n15012);
   U13546 : OAI221_X1 port map( B1 => n11742, B2 => n366, C1 => n11006, C2 => 
                           n377, A => n15026, ZN => n15025);
   U13547 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_31_15_port, B1 => 
                           n399, B2 => REGISTERS_35_15_port, C1 => n410, C2 => 
                           REGISTERS_39_15_port, ZN => n15026);
   U13548 : OAI221_X1 port map( B1 => n11582, B2 => n421, C1 => n11710, C2 => 
                           n432, A => n15027, ZN => n15024);
   U13549 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_26_15_port, B1 => 
                           n454, B2 => REGISTERS_30_15_port, C1 => n465, C2 => 
                           REGISTERS_34_15_port, ZN => n15027);
   U13550 : OAI221_X1 port map( B1 => n11422, B2 => n476, C1 => n11550, C2 => 
                           n487, A => n15028, ZN => n15023);
   U13551 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_21_15_port, B1 => 
                           n509, B2 => REGISTERS_25_15_port, C1 => n520, C2 => 
                           REGISTERS_29_15_port, ZN => n15028);
   U13552 : OAI221_X1 port map( B1 => n11262, B2 => n531, C1 => n11390, C2 => 
                           n542, A => n15029, ZN => n15022);
   U13553 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_24_15_port, B1 => 
                           n564, B2 => REGISTERS_22_15_port, C1 => n575, C2 => 
                           REGISTERS_20_15_port, ZN => n15029);
   U13554 : AOI22_X1 port map( A1 => n13880, A2 => n5024, B1 => n13881, B2 => 
                           n5025, ZN => n14990);
   U13555 : NOR4_X1 port map( A1 => n15032, A2 => n15033, A3 => n15034, A4 => 
                           n15035, ZN => n15031);
   U13556 : OAI221_X1 port map( B1 => n11070, B2 => n311, C1 => n11006, C2 => 
                           n322, A => n15036, ZN => n15035);
   U13557 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_14_15_port, B1 => 
                           n13808, B2 => REGISTERS_38_15_port, C1 => n13889, C2
                           => REGISTERS_39_15_port, ZN => n15036);
   U13558 : OAI221_X1 port map( B1 => n10910, B2 => n13810, C1 => n10846, C2 =>
                           n13890, A => n15037, ZN => n15034);
   U13559 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_15_port, B1 => 
                           n343, B2 => REGISTERS_9_15_port, C1 => n13812, C2 =>
                           REGISTERS_16_15_port, ZN => n15037);
   U13560 : OAI221_X1 port map( B1 => n10750, B2 => n303, C1 => n10686, C2 => 
                           n13893, A => n15038, ZN => n15033);
   U13561 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_15_port, B1 => 
                           n354, B2 => REGISTERS_4_15_port, C1 => n13818, C2 =>
                           REGISTERS_11_15_port, ZN => n15038);
   U13562 : OAI221_X1 port map( B1 => n11614, B2 => n304, C1 => n10558, C2 => 
                           n13896, A => n15039, ZN => n15032);
   U13563 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_15_port, B1 => 
                           n13826, B2 => REGISTERS_0_15_port, C1 => n13824, C2 
                           => REGISTERS_6_15_port, ZN => n15039);
   U13564 : NOR4_X1 port map( A1 => n15040, A2 => n15041, A3 => n15042, A4 => 
                           n15043, ZN => n15030);
   U13565 : OAI221_X1 port map( B1 => n11678, B2 => n366, C1 => n10942, C2 => 
                           n377, A => n15044, ZN => n15043);
   U13566 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_29_15_port, B1 => 
                           n399, B2 => REGISTERS_33_15_port, C1 => n410, C2 => 
                           REGISTERS_37_15_port, ZN => n15044);
   U13567 : OAI221_X1 port map( B1 => n11518, B2 => n421, C1 => n11646, C2 => 
                           n432, A => n15045, ZN => n15042);
   U13568 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_24_15_port, B1 => 
                           n454, B2 => REGISTERS_28_15_port, C1 => n465, C2 => 
                           REGISTERS_32_15_port, ZN => n15045);
   U13569 : OAI221_X1 port map( B1 => n11358, B2 => n476, C1 => n11486, C2 => 
                           n487, A => n15046, ZN => n15041);
   U13570 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_19_15_port, B1 => 
                           n509, B2 => REGISTERS_23_15_port, C1 => n520, C2 => 
                           REGISTERS_27_15_port, ZN => n15046);
   U13571 : OAI221_X1 port map( B1 => n11198, B2 => n531, C1 => n11326, C2 => 
                           n542, A => n15047, ZN => n15040);
   U13572 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_22_15_port, B1 => 
                           n564, B2 => REGISTERS_20_15_port, C1 => n575, C2 => 
                           REGISTERS_18_15_port, ZN => n15047);
   U13573 : NOR4_X1 port map( A1 => n15050, A2 => n15051, A3 => n15052, A4 => 
                           n15053, ZN => n15049);
   U13574 : OAI221_X1 port map( B1 => n11038, B2 => n311, C1 => n10974, C2 => 
                           n322, A => n15054, ZN => n15053);
   U13575 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_13_15_port, B1 => 
                           n13808, B2 => REGISTERS_37_15_port, C1 => n13889, C2
                           => REGISTERS_38_15_port, ZN => n15054);
   U13576 : OAI221_X1 port map( B1 => n10878, B2 => n13810, C1 => n10814, C2 =>
                           n13890, A => n15055, ZN => n15052);
   U13577 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_15_port, B1 => 
                           n343, B2 => REGISTERS_8_15_port, C1 => n13812, C2 =>
                           REGISTERS_15_15_port, ZN => n15055);
   U13578 : OAI221_X1 port map( B1 => n10718, B2 => n303, C1 => n10654, C2 => 
                           n13893, A => n15056, ZN => n15051);
   U13579 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_15_port, B1 => 
                           n354, B2 => REGISTERS_3_15_port, C1 => n13818, C2 =>
                           REGISTERS_10_15_port, ZN => n15056);
   U13580 : OAI221_X1 port map( B1 => n11582, B2 => n304, C1 => n10496, C2 => 
                           n13896, A => n15057, ZN => n15050);
   U13581 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_15_port, B1 => 
                           n13917, B2 => REGISTERS_39_15_port, C1 => n13824, C2
                           => REGISTERS_5_15_port, ZN => n15057);
   U13582 : NOR4_X1 port map( A1 => n15058, A2 => n15059, A3 => n15060, A4 => 
                           n15061, ZN => n15048);
   U13583 : OAI221_X1 port map( B1 => n11646, B2 => n366, C1 => n10910, C2 => 
                           n377, A => n15062, ZN => n15061);
   U13584 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_28_15_port, B1 => 
                           n399, B2 => REGISTERS_32_15_port, C1 => n410, C2 => 
                           REGISTERS_36_15_port, ZN => n15062);
   U13585 : OAI221_X1 port map( B1 => n11486, B2 => n421, C1 => n11614, C2 => 
                           n432, A => n15063, ZN => n15060);
   U13586 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_23_15_port, B1 => 
                           n454, B2 => REGISTERS_27_15_port, C1 => n465, C2 => 
                           REGISTERS_31_15_port, ZN => n15063);
   U13587 : OAI221_X1 port map( B1 => n11326, B2 => n476, C1 => n11454, C2 => 
                           n487, A => n15064, ZN => n15059);
   U13588 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_18_15_port, B1 => 
                           n509, B2 => REGISTERS_22_15_port, C1 => n520, C2 => 
                           REGISTERS_26_15_port, ZN => n15064);
   U13589 : OAI221_X1 port map( B1 => n11166, B2 => n531, C1 => n11294, C2 => 
                           n542, A => n15065, ZN => n15058);
   U13590 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_21_15_port, B1 => 
                           n564, B2 => REGISTERS_19_15_port, C1 => n575, C2 => 
                           REGISTERS_17_15_port, ZN => n15065);
   U13591 : NAND3_X1 port map( A1 => n15066, A2 => n15067, A3 => n15068, ZN => 
                           n11888);
   U13592 : AOI221_X1 port map( B1 => n13792, B2 => n5029, C1 => n13793, C2 => 
                           MEM_IN(16), A => n15069, ZN => n15068);
   U13593 : OAI22_X1 port map( A1 => n10493, A2 => n251, B1 => n5031, B2 => 
                           n121, ZN => n15069);
   U13594 : NOR2_X1 port map( A1 => n5648, A2 => n13796, ZN => n5646);
   U13595 : INV_X1 port map( A => MEM_IN(16), ZN => n5648);
   U13596 : AOI22_X1 port map( A1 => n197, A2 => n5032, B1 => n150, B2 => n5033
                           , ZN => n15067);
   U13597 : NOR4_X1 port map( A1 => n15072, A2 => n15073, A3 => n15074, A4 => 
                           n15075, ZN => n15071);
   U13598 : OAI221_X1 port map( B1 => n11101, B2 => n311, C1 => n11037, C2 => 
                           n322, A => n15076, ZN => n15075);
   U13599 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_15_16_port, B1 => 
                           n13807, B2 => REGISTERS_11_16_port, C1 => n13808, C2
                           => REGISTERS_39_16_port, ZN => n15076);
   U13600 : OAI221_X1 port map( B1 => n10813, B2 => n13809, C1 => n10941, C2 =>
                           n13810, A => n15077, ZN => n15074);
   U13601 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_16_port, B1 =>
                           n13813, B2 => REGISTERS_6_16_port, C1 => n348, C2 =>
                           REGISTERS_10_16_port, ZN => n15077);
   U13602 : OAI221_X1 port map( B1 => n10653, B2 => n13815, C1 => n10781, C2 =>
                           n303, A => n15078, ZN => n15073);
   U13603 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_16_port, B1 =>
                           n13819, B2 => REGISTERS_2_16_port, C1 => n359, C2 =>
                           REGISTERS_5_16_port, ZN => n15078);
   U13604 : OAI221_X1 port map( B1 => n10621, B2 => n13821, C1 => n11645, C2 =>
                           n304, A => n15079, ZN => n15072);
   U13605 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_16_port, B1 => 
                           n13825, B2 => REGISTERS_0_16_port, C1 => n13826, C2 
                           => REGISTERS_1_16_port, ZN => n15079);
   U13606 : NOR4_X1 port map( A1 => n15080, A2 => n15081, A3 => n15082, A4 => 
                           n15083, ZN => n15070);
   U13607 : OAI221_X1 port map( B1 => n11709, B2 => n366, C1 => n10973, C2 => 
                           n377, A => n15084, ZN => n15083);
   U13608 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_30_16_port, B1 => 
                           n399, B2 => REGISTERS_34_16_port, C1 => n410, C2 => 
                           REGISTERS_38_16_port, ZN => n15084);
   U13609 : OAI221_X1 port map( B1 => n11549, B2 => n421, C1 => n11677, C2 => 
                           n432, A => n15085, ZN => n15082);
   U13610 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_25_16_port, B1 => 
                           n454, B2 => REGISTERS_29_16_port, C1 => n465, C2 => 
                           REGISTERS_33_16_port, ZN => n15085);
   U13611 : OAI221_X1 port map( B1 => n11389, B2 => n476, C1 => n11517, C2 => 
                           n487, A => n15086, ZN => n15081);
   U13612 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_20_16_port, B1 => 
                           n509, B2 => REGISTERS_24_16_port, C1 => n520, C2 => 
                           REGISTERS_28_16_port, ZN => n15086);
   U13613 : OAI221_X1 port map( B1 => n11229, B2 => n531, C1 => n11357, C2 => 
                           n542, A => n15087, ZN => n15080);
   U13614 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_23_16_port, B1 => 
                           n564, B2 => REGISTERS_21_16_port, C1 => n575, C2 => 
                           REGISTERS_19_16_port, ZN => n15087);
   U13615 : NOR4_X1 port map( A1 => n15090, A2 => n15091, A3 => n15092, A4 => 
                           n15093, ZN => n15089);
   U13616 : OAI221_X1 port map( B1 => n11133, B2 => n311, C1 => n11069, C2 => 
                           n322, A => n15094, ZN => n15093);
   U13617 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_16_16_port, B1 => 
                           n119, B2 => REGISTERS_14_16_port, C1 => n13807, C2 
                           => REGISTERS_12_16_port, ZN => n15094);
   U13618 : OAI221_X1 port map( B1 => n11101, B2 => n13863, C1 => n10845, C2 =>
                           n13809, A => n15095, ZN => n15092);
   U13619 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_16_port, B1 => 
                           n13865, B2 => REGISTERS_9_16_port, C1 => n13813, C2 
                           => REGISTERS_7_16_port, ZN => n15095);
   U13620 : OAI221_X1 port map( B1 => n10941, B2 => n13866, C1 => n10685, C2 =>
                           n13815, A => n15096, ZN => n15091);
   U13621 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_16_port, B1 => 
                           n13868, B2 => REGISTERS_36_16_port, C1 => n13819, C2
                           => REGISTERS_3_16_port, ZN => n15096);
   U13622 : OAI221_X1 port map( B1 => n10781, B2 => n13869, C1 => n10653, C2 =>
                           n13821, A => n15097, ZN => n15090);
   U13623 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_16_port, B1 => 
                           n13871, B2 => REGISTERS_0_16_port, C1 => n13825, C2 
                           => REGISTERS_1_16_port, ZN => n15097);
   U13624 : NOR4_X1 port map( A1 => n15098, A2 => n15099, A3 => n15100, A4 => 
                           n15101, ZN => n15088);
   U13625 : OAI221_X1 port map( B1 => n11741, B2 => n366, C1 => n11005, C2 => 
                           n377, A => n15102, ZN => n15101);
   U13626 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_31_16_port, B1 => 
                           n399, B2 => REGISTERS_35_16_port, C1 => n410, C2 => 
                           REGISTERS_39_16_port, ZN => n15102);
   U13627 : OAI221_X1 port map( B1 => n11581, B2 => n421, C1 => n11709, C2 => 
                           n432, A => n15103, ZN => n15100);
   U13628 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_26_16_port, B1 => 
                           n454, B2 => REGISTERS_30_16_port, C1 => n465, C2 => 
                           REGISTERS_34_16_port, ZN => n15103);
   U13629 : OAI221_X1 port map( B1 => n11421, B2 => n476, C1 => n11549, C2 => 
                           n487, A => n15104, ZN => n15099);
   U13630 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_21_16_port, B1 => 
                           n509, B2 => REGISTERS_25_16_port, C1 => n520, C2 => 
                           REGISTERS_29_16_port, ZN => n15104);
   U13631 : OAI221_X1 port map( B1 => n11261, B2 => n531, C1 => n11389, C2 => 
                           n542, A => n15105, ZN => n15098);
   U13632 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_24_16_port, B1 => 
                           n564, B2 => REGISTERS_22_16_port, C1 => n575, C2 => 
                           REGISTERS_20_16_port, ZN => n15105);
   U13633 : AOI22_X1 port map( A1 => n13880, A2 => n5034, B1 => n13881, B2 => 
                           n5035, ZN => n15066);
   U13634 : NOR4_X1 port map( A1 => n15108, A2 => n15109, A3 => n15110, A4 => 
                           n15111, ZN => n15107);
   U13635 : OAI221_X1 port map( B1 => n11069, B2 => n311, C1 => n11005, C2 => 
                           n322, A => n15112, ZN => n15111);
   U13636 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_14_16_port, B1 => 
                           n13808, B2 => REGISTERS_38_16_port, C1 => n13889, C2
                           => REGISTERS_39_16_port, ZN => n15112);
   U13637 : OAI221_X1 port map( B1 => n10909, B2 => n13810, C1 => n10845, C2 =>
                           n13890, A => n15113, ZN => n15110);
   U13638 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_16_port, B1 => 
                           n343, B2 => REGISTERS_9_16_port, C1 => n13812, C2 =>
                           REGISTERS_16_16_port, ZN => n15113);
   U13639 : OAI221_X1 port map( B1 => n10749, B2 => n303, C1 => n10685, C2 => 
                           n13893, A => n15114, ZN => n15109);
   U13640 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_16_port, B1 => 
                           n354, B2 => REGISTERS_4_16_port, C1 => n13818, C2 =>
                           REGISTERS_11_16_port, ZN => n15114);
   U13641 : OAI221_X1 port map( B1 => n11613, B2 => n304, C1 => n10557, C2 => 
                           n13896, A => n15115, ZN => n15108);
   U13642 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_16_port, B1 => 
                           n13826, B2 => REGISTERS_0_16_port, C1 => n13824, C2 
                           => REGISTERS_6_16_port, ZN => n15115);
   U13643 : NOR4_X1 port map( A1 => n15116, A2 => n15117, A3 => n15118, A4 => 
                           n15119, ZN => n15106);
   U13644 : OAI221_X1 port map( B1 => n11677, B2 => n366, C1 => n10941, C2 => 
                           n377, A => n15120, ZN => n15119);
   U13645 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_29_16_port, B1 => 
                           n399, B2 => REGISTERS_33_16_port, C1 => n410, C2 => 
                           REGISTERS_37_16_port, ZN => n15120);
   U13646 : OAI221_X1 port map( B1 => n11517, B2 => n421, C1 => n11645, C2 => 
                           n432, A => n15121, ZN => n15118);
   U13647 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_24_16_port, B1 => 
                           n454, B2 => REGISTERS_28_16_port, C1 => n465, C2 => 
                           REGISTERS_32_16_port, ZN => n15121);
   U13648 : OAI221_X1 port map( B1 => n11357, B2 => n476, C1 => n11485, C2 => 
                           n487, A => n15122, ZN => n15117);
   U13649 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_19_16_port, B1 => 
                           n509, B2 => REGISTERS_23_16_port, C1 => n520, C2 => 
                           REGISTERS_27_16_port, ZN => n15122);
   U13650 : OAI221_X1 port map( B1 => n11197, B2 => n531, C1 => n11325, C2 => 
                           n542, A => n15123, ZN => n15116);
   U13651 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_22_16_port, B1 => 
                           n564, B2 => REGISTERS_20_16_port, C1 => n575, C2 => 
                           REGISTERS_18_16_port, ZN => n15123);
   U13652 : NOR4_X1 port map( A1 => n15126, A2 => n15127, A3 => n15128, A4 => 
                           n15129, ZN => n15125);
   U13653 : OAI221_X1 port map( B1 => n11037, B2 => n311, C1 => n10973, C2 => 
                           n322, A => n15130, ZN => n15129);
   U13654 : AOI222_X1 port map( A1 => n333, A2 => REGISTERS_13_16_port, B1 => 
                           n13808, B2 => REGISTERS_37_16_port, C1 => n13889, C2
                           => REGISTERS_38_16_port, ZN => n15130);
   U13655 : OAI221_X1 port map( B1 => n10877, B2 => n13810, C1 => n10813, C2 =>
                           n13890, A => n15131, ZN => n15128);
   U13656 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_16_port, B1 => 
                           n343, B2 => REGISTERS_8_16_port, C1 => n13812, C2 =>
                           REGISTERS_15_16_port, ZN => n15131);
   U13657 : OAI221_X1 port map( B1 => n10717, B2 => n303, C1 => n10653, C2 => 
                           n13893, A => n15132, ZN => n15127);
   U13658 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_16_port, B1 => 
                           n354, B2 => REGISTERS_3_16_port, C1 => n13818, C2 =>
                           REGISTERS_10_16_port, ZN => n15132);
   U13659 : OAI221_X1 port map( B1 => n11581, B2 => n304, C1 => n10493, C2 => 
                           n13896, A => n15133, ZN => n15126);
   U13660 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_16_port, B1 => 
                           n13917, B2 => REGISTERS_39_16_port, C1 => n13824, C2
                           => REGISTERS_5_16_port, ZN => n15133);
   U13661 : NOR4_X1 port map( A1 => n15134, A2 => n15135, A3 => n15136, A4 => 
                           n15137, ZN => n15124);
   U13662 : OAI221_X1 port map( B1 => n11645, B2 => n366, C1 => n10909, C2 => 
                           n377, A => n15138, ZN => n15137);
   U13663 : AOI222_X1 port map( A1 => n388, A2 => REGISTERS_28_16_port, B1 => 
                           n399, B2 => REGISTERS_32_16_port, C1 => n410, C2 => 
                           REGISTERS_36_16_port, ZN => n15138);
   U13664 : OAI221_X1 port map( B1 => n11485, B2 => n421, C1 => n11613, C2 => 
                           n432, A => n15139, ZN => n15136);
   U13665 : AOI222_X1 port map( A1 => n443, A2 => REGISTERS_23_16_port, B1 => 
                           n454, B2 => REGISTERS_27_16_port, C1 => n465, C2 => 
                           REGISTERS_31_16_port, ZN => n15139);
   U13666 : OAI221_X1 port map( B1 => n11325, B2 => n476, C1 => n11453, C2 => 
                           n487, A => n15140, ZN => n15135);
   U13667 : AOI222_X1 port map( A1 => n498, A2 => REGISTERS_18_16_port, B1 => 
                           n509, B2 => REGISTERS_22_16_port, C1 => n520, C2 => 
                           REGISTERS_26_16_port, ZN => n15140);
   U13668 : OAI221_X1 port map( B1 => n11165, B2 => n531, C1 => n11293, C2 => 
                           n542, A => n15141, ZN => n15134);
   U13669 : AOI222_X1 port map( A1 => n553, A2 => REGISTERS_21_16_port, B1 => 
                           n564, B2 => REGISTERS_19_16_port, C1 => n575, C2 => 
                           REGISTERS_17_16_port, ZN => n15141);
   U13670 : NAND3_X1 port map( A1 => n15142, A2 => n15143, A3 => n15144, ZN => 
                           n11887);
   U13671 : AOI221_X1 port map( B1 => n13792, B2 => n5039, C1 => n13793, C2 => 
                           MEM_IN(17), A => n15145, ZN => n15144);
   U13672 : OAI22_X1 port map( A1 => n10490, A2 => n251, B1 => n5041, B2 => 
                           n121, ZN => n15145);
   U13673 : NOR2_X1 port map( A1 => n5655, A2 => n13796, ZN => n5653);
   U13674 : INV_X1 port map( A => MEM_IN(17), ZN => n5655);
   U13675 : AOI22_X1 port map( A1 => n197, A2 => n5042, B1 => n150, B2 => n5043
                           , ZN => n15143);
   U13676 : NOR4_X1 port map( A1 => n15148, A2 => n15149, A3 => n15150, A4 => 
                           n15151, ZN => n15147);
   U13677 : OAI221_X1 port map( B1 => n11100, B2 => n310, C1 => n11036, C2 => 
                           n321, A => n15152, ZN => n15151);
   U13678 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_15_17_port, B1 => 
                           n13807, B2 => REGISTERS_11_17_port, C1 => n13808, C2
                           => REGISTERS_39_17_port, ZN => n15152);
   U13679 : OAI221_X1 port map( B1 => n10812, B2 => n13809, C1 => n10940, C2 =>
                           n13810, A => n15153, ZN => n15150);
   U13680 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_17_port, B1 =>
                           n13813, B2 => REGISTERS_6_17_port, C1 => n348, C2 =>
                           REGISTERS_10_17_port, ZN => n15153);
   U13681 : OAI221_X1 port map( B1 => n10652, B2 => n13815, C1 => n10780, C2 =>
                           n303, A => n15154, ZN => n15149);
   U13682 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_17_port, B1 =>
                           n13819, B2 => REGISTERS_2_17_port, C1 => n359, C2 =>
                           REGISTERS_5_17_port, ZN => n15154);
   U13683 : OAI221_X1 port map( B1 => n10620, B2 => n13821, C1 => n11644, C2 =>
                           n304, A => n15155, ZN => n15148);
   U13684 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_17_port, B1 => 
                           n13825, B2 => REGISTERS_0_17_port, C1 => n13826, C2 
                           => REGISTERS_1_17_port, ZN => n15155);
   U13685 : NOR4_X1 port map( A1 => n15156, A2 => n15157, A3 => n15158, A4 => 
                           n15159, ZN => n15146);
   U13686 : OAI221_X1 port map( B1 => n11708, B2 => n365, C1 => n10972, C2 => 
                           n377, A => n15160, ZN => n15159);
   U13687 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_30_17_port, B1 => 
                           n398, B2 => REGISTERS_34_17_port, C1 => n409, C2 => 
                           REGISTERS_38_17_port, ZN => n15160);
   U13688 : OAI221_X1 port map( B1 => n11548, B2 => n420, C1 => n11676, C2 => 
                           n431, A => n15161, ZN => n15158);
   U13689 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_25_17_port, B1 => 
                           n453, B2 => REGISTERS_29_17_port, C1 => n464, C2 => 
                           REGISTERS_33_17_port, ZN => n15161);
   U13690 : OAI221_X1 port map( B1 => n11388, B2 => n475, C1 => n11516, C2 => 
                           n486, A => n15162, ZN => n15157);
   U13691 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_20_17_port, B1 => 
                           n508, B2 => REGISTERS_24_17_port, C1 => n519, C2 => 
                           REGISTERS_28_17_port, ZN => n15162);
   U13692 : OAI221_X1 port map( B1 => n11228, B2 => n530, C1 => n11356, C2 => 
                           n541, A => n15163, ZN => n15156);
   U13693 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_23_17_port, B1 => 
                           n563, B2 => REGISTERS_21_17_port, C1 => n574, C2 => 
                           REGISTERS_19_17_port, ZN => n15163);
   U13694 : NOR4_X1 port map( A1 => n15166, A2 => n15167, A3 => n15168, A4 => 
                           n15169, ZN => n15165);
   U13695 : OAI221_X1 port map( B1 => n11132, B2 => n310, C1 => n11068, C2 => 
                           n321, A => n15170, ZN => n15169);
   U13696 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_16_17_port, B1 => 
                           n119, B2 => REGISTERS_14_17_port, C1 => n13807, C2 
                           => REGISTERS_12_17_port, ZN => n15170);
   U13697 : OAI221_X1 port map( B1 => n11100, B2 => n13863, C1 => n10844, C2 =>
                           n13809, A => n15171, ZN => n15168);
   U13698 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_17_port, B1 => 
                           n13865, B2 => REGISTERS_9_17_port, C1 => n13813, C2 
                           => REGISTERS_7_17_port, ZN => n15171);
   U13699 : OAI221_X1 port map( B1 => n10940, B2 => n13866, C1 => n10684, C2 =>
                           n13815, A => n15172, ZN => n15167);
   U13700 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_17_port, B1 => 
                           n13868, B2 => REGISTERS_36_17_port, C1 => n13819, C2
                           => REGISTERS_3_17_port, ZN => n15172);
   U13701 : OAI221_X1 port map( B1 => n10780, B2 => n13869, C1 => n10652, C2 =>
                           n13821, A => n15173, ZN => n15166);
   U13702 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_17_port, B1 => 
                           n13871, B2 => REGISTERS_0_17_port, C1 => n13825, C2 
                           => REGISTERS_1_17_port, ZN => n15173);
   U13703 : NOR4_X1 port map( A1 => n15174, A2 => n15175, A3 => n15176, A4 => 
                           n15177, ZN => n15164);
   U13704 : OAI221_X1 port map( B1 => n11740, B2 => n365, C1 => n11004, C2 => 
                           n376, A => n15178, ZN => n15177);
   U13705 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_31_17_port, B1 => 
                           n398, B2 => REGISTERS_35_17_port, C1 => n409, C2 => 
                           REGISTERS_39_17_port, ZN => n15178);
   U13706 : OAI221_X1 port map( B1 => n11580, B2 => n420, C1 => n11708, C2 => 
                           n431, A => n15179, ZN => n15176);
   U13707 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_26_17_port, B1 => 
                           n453, B2 => REGISTERS_30_17_port, C1 => n464, C2 => 
                           REGISTERS_34_17_port, ZN => n15179);
   U13708 : OAI221_X1 port map( B1 => n11420, B2 => n475, C1 => n11548, C2 => 
                           n486, A => n15180, ZN => n15175);
   U13709 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_21_17_port, B1 => 
                           n508, B2 => REGISTERS_25_17_port, C1 => n519, C2 => 
                           REGISTERS_29_17_port, ZN => n15180);
   U13710 : OAI221_X1 port map( B1 => n11260, B2 => n530, C1 => n11388, C2 => 
                           n541, A => n15181, ZN => n15174);
   U13711 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_24_17_port, B1 => 
                           n563, B2 => REGISTERS_22_17_port, C1 => n574, C2 => 
                           REGISTERS_20_17_port, ZN => n15181);
   U13712 : AOI22_X1 port map( A1 => n13880, A2 => n5044, B1 => n13881, B2 => 
                           n5045, ZN => n15142);
   U13713 : NOR4_X1 port map( A1 => n15184, A2 => n15185, A3 => n15186, A4 => 
                           n15187, ZN => n15183);
   U13714 : OAI221_X1 port map( B1 => n11068, B2 => n310, C1 => n11004, C2 => 
                           n321, A => n15188, ZN => n15187);
   U13715 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_14_17_port, B1 => 
                           n13808, B2 => REGISTERS_38_17_port, C1 => n13889, C2
                           => REGISTERS_39_17_port, ZN => n15188);
   U13716 : OAI221_X1 port map( B1 => n10908, B2 => n13810, C1 => n10844, C2 =>
                           n13890, A => n15189, ZN => n15186);
   U13717 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_17_port, B1 => 
                           n344, B2 => REGISTERS_9_17_port, C1 => n13812, C2 =>
                           REGISTERS_16_17_port, ZN => n15189);
   U13718 : OAI221_X1 port map( B1 => n10748, B2 => n303, C1 => n10684, C2 => 
                           n13893, A => n15190, ZN => n15185);
   U13719 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_17_port, B1 => 
                           n355, B2 => REGISTERS_4_17_port, C1 => n13818, C2 =>
                           REGISTERS_11_17_port, ZN => n15190);
   U13720 : OAI221_X1 port map( B1 => n11612, B2 => n304, C1 => n10556, C2 => 
                           n13896, A => n15191, ZN => n15184);
   U13721 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_17_port, B1 => 
                           n13826, B2 => REGISTERS_0_17_port, C1 => n13824, C2 
                           => REGISTERS_6_17_port, ZN => n15191);
   U13722 : NOR4_X1 port map( A1 => n15192, A2 => n15193, A3 => n15194, A4 => 
                           n15195, ZN => n15182);
   U13723 : OAI221_X1 port map( B1 => n11676, B2 => n365, C1 => n10940, C2 => 
                           n376, A => n15196, ZN => n15195);
   U13724 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_29_17_port, B1 => 
                           n398, B2 => REGISTERS_33_17_port, C1 => n409, C2 => 
                           REGISTERS_37_17_port, ZN => n15196);
   U13725 : OAI221_X1 port map( B1 => n11516, B2 => n420, C1 => n11644, C2 => 
                           n431, A => n15197, ZN => n15194);
   U13726 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_24_17_port, B1 => 
                           n453, B2 => REGISTERS_28_17_port, C1 => n464, C2 => 
                           REGISTERS_32_17_port, ZN => n15197);
   U13727 : OAI221_X1 port map( B1 => n11356, B2 => n475, C1 => n11484, C2 => 
                           n486, A => n15198, ZN => n15193);
   U13728 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_19_17_port, B1 => 
                           n508, B2 => REGISTERS_23_17_port, C1 => n519, C2 => 
                           REGISTERS_27_17_port, ZN => n15198);
   U13729 : OAI221_X1 port map( B1 => n11196, B2 => n530, C1 => n11324, C2 => 
                           n541, A => n15199, ZN => n15192);
   U13730 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_22_17_port, B1 => 
                           n563, B2 => REGISTERS_20_17_port, C1 => n574, C2 => 
                           REGISTERS_18_17_port, ZN => n15199);
   U13731 : NOR4_X1 port map( A1 => n15202, A2 => n15203, A3 => n15204, A4 => 
                           n15205, ZN => n15201);
   U13732 : OAI221_X1 port map( B1 => n11036, B2 => n310, C1 => n10972, C2 => 
                           n321, A => n15206, ZN => n15205);
   U13733 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_13_17_port, B1 => 
                           n13808, B2 => REGISTERS_37_17_port, C1 => n13889, C2
                           => REGISTERS_38_17_port, ZN => n15206);
   U13734 : OAI221_X1 port map( B1 => n10876, B2 => n13810, C1 => n10812, C2 =>
                           n13890, A => n15207, ZN => n15204);
   U13735 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_17_port, B1 => 
                           n344, B2 => REGISTERS_8_17_port, C1 => n13812, C2 =>
                           REGISTERS_15_17_port, ZN => n15207);
   U13736 : OAI221_X1 port map( B1 => n10716, B2 => n303, C1 => n10652, C2 => 
                           n13893, A => n15208, ZN => n15203);
   U13737 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_17_port, B1 => 
                           n355, B2 => REGISTERS_3_17_port, C1 => n13818, C2 =>
                           REGISTERS_10_17_port, ZN => n15208);
   U13738 : OAI221_X1 port map( B1 => n11580, B2 => n304, C1 => n10490, C2 => 
                           n13896, A => n15209, ZN => n15202);
   U13739 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_17_port, B1 => 
                           n13917, B2 => REGISTERS_39_17_port, C1 => n13824, C2
                           => REGISTERS_5_17_port, ZN => n15209);
   U13740 : NOR4_X1 port map( A1 => n15210, A2 => n15211, A3 => n15212, A4 => 
                           n15213, ZN => n15200);
   U13741 : OAI221_X1 port map( B1 => n11644, B2 => n365, C1 => n10908, C2 => 
                           n376, A => n15214, ZN => n15213);
   U13742 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_28_17_port, B1 => 
                           n398, B2 => REGISTERS_32_17_port, C1 => n409, C2 => 
                           REGISTERS_36_17_port, ZN => n15214);
   U13743 : OAI221_X1 port map( B1 => n11484, B2 => n420, C1 => n11612, C2 => 
                           n431, A => n15215, ZN => n15212);
   U13744 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_23_17_port, B1 => 
                           n453, B2 => REGISTERS_27_17_port, C1 => n464, C2 => 
                           REGISTERS_31_17_port, ZN => n15215);
   U13745 : OAI221_X1 port map( B1 => n11324, B2 => n475, C1 => n11452, C2 => 
                           n486, A => n15216, ZN => n15211);
   U13746 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_18_17_port, B1 => 
                           n508, B2 => REGISTERS_22_17_port, C1 => n519, C2 => 
                           REGISTERS_26_17_port, ZN => n15216);
   U13747 : OAI221_X1 port map( B1 => n11164, B2 => n530, C1 => n11292, C2 => 
                           n541, A => n15217, ZN => n15210);
   U13748 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_21_17_port, B1 => 
                           n563, B2 => REGISTERS_19_17_port, C1 => n574, C2 => 
                           REGISTERS_17_17_port, ZN => n15217);
   U13749 : NAND3_X1 port map( A1 => n15218, A2 => n15219, A3 => n15220, ZN => 
                           n11886);
   U13750 : AOI221_X1 port map( B1 => n13792, B2 => n5049, C1 => n13793, C2 => 
                           MEM_IN(18), A => n15221, ZN => n15220);
   U13751 : OAI22_X1 port map( A1 => n10487, A2 => n251, B1 => n5051, B2 => 
                           n121, ZN => n15221);
   U13752 : NOR2_X1 port map( A1 => n5662, A2 => n13796, ZN => n5660);
   U13753 : INV_X1 port map( A => MEM_IN(18), ZN => n5662);
   U13754 : AOI22_X1 port map( A1 => n197, A2 => n5052, B1 => n150, B2 => n5053
                           , ZN => n15219);
   U13755 : NOR4_X1 port map( A1 => n15224, A2 => n15225, A3 => n15226, A4 => 
                           n15227, ZN => n15223);
   U13756 : OAI221_X1 port map( B1 => n11099, B2 => n310, C1 => n11035, C2 => 
                           n321, A => n15228, ZN => n15227);
   U13757 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_15_18_port, B1 => 
                           n13807, B2 => REGISTERS_11_18_port, C1 => n13808, C2
                           => REGISTERS_39_18_port, ZN => n15228);
   U13758 : OAI221_X1 port map( B1 => n10811, B2 => n13809, C1 => n10939, C2 =>
                           n13810, A => n15229, ZN => n15226);
   U13759 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_18_port, B1 =>
                           n13813, B2 => REGISTERS_6_18_port, C1 => n348, C2 =>
                           REGISTERS_10_18_port, ZN => n15229);
   U13760 : OAI221_X1 port map( B1 => n10651, B2 => n13815, C1 => n10779, C2 =>
                           n303, A => n15230, ZN => n15225);
   U13761 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_18_port, B1 =>
                           n13819, B2 => REGISTERS_2_18_port, C1 => n359, C2 =>
                           REGISTERS_5_18_port, ZN => n15230);
   U13762 : OAI221_X1 port map( B1 => n10619, B2 => n13821, C1 => n11643, C2 =>
                           n304, A => n15231, ZN => n15224);
   U13763 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_18_port, B1 => 
                           n13825, B2 => REGISTERS_0_18_port, C1 => n13826, C2 
                           => REGISTERS_1_18_port, ZN => n15231);
   U13764 : NOR4_X1 port map( A1 => n15232, A2 => n15233, A3 => n15234, A4 => 
                           n15235, ZN => n15222);
   U13765 : OAI221_X1 port map( B1 => n11707, B2 => n365, C1 => n10971, C2 => 
                           n376, A => n15236, ZN => n15235);
   U13766 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_30_18_port, B1 => 
                           n398, B2 => REGISTERS_34_18_port, C1 => n409, C2 => 
                           REGISTERS_38_18_port, ZN => n15236);
   U13767 : OAI221_X1 port map( B1 => n11547, B2 => n420, C1 => n11675, C2 => 
                           n431, A => n15237, ZN => n15234);
   U13768 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_25_18_port, B1 => 
                           n453, B2 => REGISTERS_29_18_port, C1 => n464, C2 => 
                           REGISTERS_33_18_port, ZN => n15237);
   U13769 : OAI221_X1 port map( B1 => n11387, B2 => n475, C1 => n11515, C2 => 
                           n486, A => n15238, ZN => n15233);
   U13770 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_20_18_port, B1 => 
                           n508, B2 => REGISTERS_24_18_port, C1 => n519, C2 => 
                           REGISTERS_28_18_port, ZN => n15238);
   U13771 : OAI221_X1 port map( B1 => n11227, B2 => n530, C1 => n11355, C2 => 
                           n541, A => n15239, ZN => n15232);
   U13772 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_23_18_port, B1 => 
                           n563, B2 => REGISTERS_21_18_port, C1 => n574, C2 => 
                           REGISTERS_19_18_port, ZN => n15239);
   U13773 : NOR4_X1 port map( A1 => n15242, A2 => n15243, A3 => n15244, A4 => 
                           n15245, ZN => n15241);
   U13774 : OAI221_X1 port map( B1 => n11131, B2 => n310, C1 => n11067, C2 => 
                           n321, A => n15246, ZN => n15245);
   U13775 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_16_18_port, B1 => 
                           n119, B2 => REGISTERS_14_18_port, C1 => n13807, C2 
                           => REGISTERS_12_18_port, ZN => n15246);
   U13776 : OAI221_X1 port map( B1 => n11099, B2 => n13863, C1 => n10843, C2 =>
                           n13809, A => n15247, ZN => n15244);
   U13777 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_18_port, B1 => 
                           n13865, B2 => REGISTERS_9_18_port, C1 => n13813, C2 
                           => REGISTERS_7_18_port, ZN => n15247);
   U13778 : OAI221_X1 port map( B1 => n10939, B2 => n13866, C1 => n10683, C2 =>
                           n13815, A => n15248, ZN => n15243);
   U13779 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_18_port, B1 => 
                           n13868, B2 => REGISTERS_36_18_port, C1 => n13819, C2
                           => REGISTERS_3_18_port, ZN => n15248);
   U13780 : OAI221_X1 port map( B1 => n10779, B2 => n13869, C1 => n10651, C2 =>
                           n13821, A => n15249, ZN => n15242);
   U13781 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_18_port, B1 => 
                           n13871, B2 => REGISTERS_0_18_port, C1 => n13825, C2 
                           => REGISTERS_1_18_port, ZN => n15249);
   U13782 : NOR4_X1 port map( A1 => n15250, A2 => n15251, A3 => n15252, A4 => 
                           n15253, ZN => n15240);
   U13783 : OAI221_X1 port map( B1 => n11739, B2 => n365, C1 => n11003, C2 => 
                           n376, A => n15254, ZN => n15253);
   U13784 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_31_18_port, B1 => 
                           n398, B2 => REGISTERS_35_18_port, C1 => n409, C2 => 
                           REGISTERS_39_18_port, ZN => n15254);
   U13785 : OAI221_X1 port map( B1 => n11579, B2 => n420, C1 => n11707, C2 => 
                           n431, A => n15255, ZN => n15252);
   U13786 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_26_18_port, B1 => 
                           n453, B2 => REGISTERS_30_18_port, C1 => n464, C2 => 
                           REGISTERS_34_18_port, ZN => n15255);
   U13787 : OAI221_X1 port map( B1 => n11419, B2 => n475, C1 => n11547, C2 => 
                           n486, A => n15256, ZN => n15251);
   U13788 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_21_18_port, B1 => 
                           n508, B2 => REGISTERS_25_18_port, C1 => n519, C2 => 
                           REGISTERS_29_18_port, ZN => n15256);
   U13789 : OAI221_X1 port map( B1 => n11259, B2 => n530, C1 => n11387, C2 => 
                           n541, A => n15257, ZN => n15250);
   U13790 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_24_18_port, B1 => 
                           n563, B2 => REGISTERS_22_18_port, C1 => n574, C2 => 
                           REGISTERS_20_18_port, ZN => n15257);
   U13791 : AOI22_X1 port map( A1 => n13880, A2 => n5054, B1 => n13881, B2 => 
                           n5055, ZN => n15218);
   U13792 : NOR4_X1 port map( A1 => n15260, A2 => n15261, A3 => n15262, A4 => 
                           n15263, ZN => n15259);
   U13793 : OAI221_X1 port map( B1 => n11067, B2 => n310, C1 => n11003, C2 => 
                           n321, A => n15264, ZN => n15263);
   U13794 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_14_18_port, B1 => 
                           n13808, B2 => REGISTERS_38_18_port, C1 => n13889, C2
                           => REGISTERS_39_18_port, ZN => n15264);
   U13795 : OAI221_X1 port map( B1 => n10907, B2 => n13810, C1 => n10843, C2 =>
                           n13890, A => n15265, ZN => n15262);
   U13796 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_18_port, B1 => 
                           n344, B2 => REGISTERS_9_18_port, C1 => n13812, C2 =>
                           REGISTERS_16_18_port, ZN => n15265);
   U13797 : OAI221_X1 port map( B1 => n10747, B2 => n303, C1 => n10683, C2 => 
                           n13893, A => n15266, ZN => n15261);
   U13798 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_18_port, B1 => 
                           n355, B2 => REGISTERS_4_18_port, C1 => n13818, C2 =>
                           REGISTERS_11_18_port, ZN => n15266);
   U13799 : OAI221_X1 port map( B1 => n11611, B2 => n304, C1 => n10555, C2 => 
                           n13896, A => n15267, ZN => n15260);
   U13800 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_18_port, B1 => 
                           n13826, B2 => REGISTERS_0_18_port, C1 => n13824, C2 
                           => REGISTERS_6_18_port, ZN => n15267);
   U13801 : NOR4_X1 port map( A1 => n15268, A2 => n15269, A3 => n15270, A4 => 
                           n15271, ZN => n15258);
   U13802 : OAI221_X1 port map( B1 => n11675, B2 => n365, C1 => n10939, C2 => 
                           n376, A => n15272, ZN => n15271);
   U13803 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_29_18_port, B1 => 
                           n398, B2 => REGISTERS_33_18_port, C1 => n409, C2 => 
                           REGISTERS_37_18_port, ZN => n15272);
   U13804 : OAI221_X1 port map( B1 => n11515, B2 => n420, C1 => n11643, C2 => 
                           n431, A => n15273, ZN => n15270);
   U13805 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_24_18_port, B1 => 
                           n453, B2 => REGISTERS_28_18_port, C1 => n464, C2 => 
                           REGISTERS_32_18_port, ZN => n15273);
   U13806 : OAI221_X1 port map( B1 => n11355, B2 => n475, C1 => n11483, C2 => 
                           n486, A => n15274, ZN => n15269);
   U13807 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_19_18_port, B1 => 
                           n508, B2 => REGISTERS_23_18_port, C1 => n519, C2 => 
                           REGISTERS_27_18_port, ZN => n15274);
   U13808 : OAI221_X1 port map( B1 => n11195, B2 => n530, C1 => n11323, C2 => 
                           n541, A => n15275, ZN => n15268);
   U13809 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_22_18_port, B1 => 
                           n563, B2 => REGISTERS_20_18_port, C1 => n574, C2 => 
                           REGISTERS_18_18_port, ZN => n15275);
   U13810 : NOR4_X1 port map( A1 => n15278, A2 => n15279, A3 => n15280, A4 => 
                           n15281, ZN => n15277);
   U13811 : OAI221_X1 port map( B1 => n11035, B2 => n310, C1 => n10971, C2 => 
                           n321, A => n15282, ZN => n15281);
   U13812 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_13_18_port, B1 => 
                           n13808, B2 => REGISTERS_37_18_port, C1 => n13889, C2
                           => REGISTERS_38_18_port, ZN => n15282);
   U13813 : OAI221_X1 port map( B1 => n10875, B2 => n13810, C1 => n10811, C2 =>
                           n13890, A => n15283, ZN => n15280);
   U13814 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_18_port, B1 => 
                           n344, B2 => REGISTERS_8_18_port, C1 => n13812, C2 =>
                           REGISTERS_15_18_port, ZN => n15283);
   U13815 : OAI221_X1 port map( B1 => n10715, B2 => n303, C1 => n10651, C2 => 
                           n13893, A => n15284, ZN => n15279);
   U13816 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_18_port, B1 => 
                           n355, B2 => REGISTERS_3_18_port, C1 => n13818, C2 =>
                           REGISTERS_10_18_port, ZN => n15284);
   U13817 : OAI221_X1 port map( B1 => n11579, B2 => n304, C1 => n10487, C2 => 
                           n13896, A => n15285, ZN => n15278);
   U13818 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_18_port, B1 => 
                           n13917, B2 => REGISTERS_39_18_port, C1 => n13824, C2
                           => REGISTERS_5_18_port, ZN => n15285);
   U13819 : NOR4_X1 port map( A1 => n15286, A2 => n15287, A3 => n15288, A4 => 
                           n15289, ZN => n15276);
   U13820 : OAI221_X1 port map( B1 => n11643, B2 => n365, C1 => n10907, C2 => 
                           n376, A => n15290, ZN => n15289);
   U13821 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_28_18_port, B1 => 
                           n398, B2 => REGISTERS_32_18_port, C1 => n409, C2 => 
                           REGISTERS_36_18_port, ZN => n15290);
   U13822 : OAI221_X1 port map( B1 => n11483, B2 => n420, C1 => n11611, C2 => 
                           n431, A => n15291, ZN => n15288);
   U13823 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_23_18_port, B1 => 
                           n453, B2 => REGISTERS_27_18_port, C1 => n464, C2 => 
                           REGISTERS_31_18_port, ZN => n15291);
   U13824 : OAI221_X1 port map( B1 => n11323, B2 => n475, C1 => n11451, C2 => 
                           n486, A => n15292, ZN => n15287);
   U13825 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_18_18_port, B1 => 
                           n508, B2 => REGISTERS_22_18_port, C1 => n519, C2 => 
                           REGISTERS_26_18_port, ZN => n15292);
   U13826 : OAI221_X1 port map( B1 => n11163, B2 => n530, C1 => n11291, C2 => 
                           n541, A => n15293, ZN => n15286);
   U13827 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_21_18_port, B1 => 
                           n563, B2 => REGISTERS_19_18_port, C1 => n574, C2 => 
                           REGISTERS_17_18_port, ZN => n15293);
   U13828 : NAND3_X1 port map( A1 => n15294, A2 => n15295, A3 => n15296, ZN => 
                           n11885);
   U13829 : AOI221_X1 port map( B1 => n13792, B2 => n5059, C1 => n13793, C2 => 
                           MEM_IN(19), A => n15297, ZN => n15296);
   U13830 : OAI22_X1 port map( A1 => n10484, A2 => n251, B1 => n5061, B2 => 
                           n121, ZN => n15297);
   U13831 : NOR2_X1 port map( A1 => n5669, A2 => n13796, ZN => n5667);
   U13832 : INV_X1 port map( A => MEM_IN(19), ZN => n5669);
   U13833 : AOI22_X1 port map( A1 => n197, A2 => n5062, B1 => n150, B2 => n5063
                           , ZN => n15295);
   U13834 : NOR4_X1 port map( A1 => n15300, A2 => n15301, A3 => n15302, A4 => 
                           n15303, ZN => n15299);
   U13835 : OAI221_X1 port map( B1 => n11098, B2 => n310, C1 => n11034, C2 => 
                           n321, A => n15304, ZN => n15303);
   U13836 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_15_19_port, B1 => 
                           n13807, B2 => REGISTERS_11_19_port, C1 => n13808, C2
                           => REGISTERS_39_19_port, ZN => n15304);
   U13837 : OAI221_X1 port map( B1 => n10810, B2 => n13809, C1 => n10938, C2 =>
                           n13810, A => n15305, ZN => n15302);
   U13838 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_19_port, B1 =>
                           n13813, B2 => REGISTERS_6_19_port, C1 => n348, C2 =>
                           REGISTERS_10_19_port, ZN => n15305);
   U13839 : OAI221_X1 port map( B1 => n10650, B2 => n13815, C1 => n10778, C2 =>
                           n303, A => n15306, ZN => n15301);
   U13840 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_19_port, B1 =>
                           n13819, B2 => REGISTERS_2_19_port, C1 => n359, C2 =>
                           REGISTERS_5_19_port, ZN => n15306);
   U13841 : OAI221_X1 port map( B1 => n10618, B2 => n13821, C1 => n11642, C2 =>
                           n304, A => n15307, ZN => n15300);
   U13842 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_19_port, B1 => 
                           n13825, B2 => REGISTERS_0_19_port, C1 => n13826, C2 
                           => REGISTERS_1_19_port, ZN => n15307);
   U13843 : NOR4_X1 port map( A1 => n15308, A2 => n15309, A3 => n15310, A4 => 
                           n15311, ZN => n15298);
   U13844 : OAI221_X1 port map( B1 => n11706, B2 => n365, C1 => n10970, C2 => 
                           n376, A => n15312, ZN => n15311);
   U13845 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_30_19_port, B1 => 
                           n398, B2 => REGISTERS_34_19_port, C1 => n409, C2 => 
                           REGISTERS_38_19_port, ZN => n15312);
   U13846 : OAI221_X1 port map( B1 => n11546, B2 => n420, C1 => n11674, C2 => 
                           n431, A => n15313, ZN => n15310);
   U13847 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_25_19_port, B1 => 
                           n453, B2 => REGISTERS_29_19_port, C1 => n464, C2 => 
                           REGISTERS_33_19_port, ZN => n15313);
   U13848 : OAI221_X1 port map( B1 => n11386, B2 => n475, C1 => n11514, C2 => 
                           n486, A => n15314, ZN => n15309);
   U13849 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_20_19_port, B1 => 
                           n508, B2 => REGISTERS_24_19_port, C1 => n519, C2 => 
                           REGISTERS_28_19_port, ZN => n15314);
   U13850 : OAI221_X1 port map( B1 => n11226, B2 => n530, C1 => n11354, C2 => 
                           n541, A => n15315, ZN => n15308);
   U13851 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_23_19_port, B1 => 
                           n563, B2 => REGISTERS_21_19_port, C1 => n574, C2 => 
                           REGISTERS_19_19_port, ZN => n15315);
   U13852 : NOR4_X1 port map( A1 => n15318, A2 => n15319, A3 => n15320, A4 => 
                           n15321, ZN => n15317);
   U13853 : OAI221_X1 port map( B1 => n11130, B2 => n310, C1 => n11066, C2 => 
                           n321, A => n15322, ZN => n15321);
   U13854 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_16_19_port, B1 => 
                           n119, B2 => REGISTERS_14_19_port, C1 => n13807, C2 
                           => REGISTERS_12_19_port, ZN => n15322);
   U13855 : OAI221_X1 port map( B1 => n11098, B2 => n13863, C1 => n10842, C2 =>
                           n13809, A => n15323, ZN => n15320);
   U13856 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_19_port, B1 => 
                           n13865, B2 => REGISTERS_9_19_port, C1 => n13813, C2 
                           => REGISTERS_7_19_port, ZN => n15323);
   U13857 : OAI221_X1 port map( B1 => n10938, B2 => n13866, C1 => n10682, C2 =>
                           n13815, A => n15324, ZN => n15319);
   U13858 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_19_port, B1 => 
                           n13868, B2 => REGISTERS_36_19_port, C1 => n13819, C2
                           => REGISTERS_3_19_port, ZN => n15324);
   U13859 : OAI221_X1 port map( B1 => n10778, B2 => n13869, C1 => n10650, C2 =>
                           n13821, A => n15325, ZN => n15318);
   U13860 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_19_port, B1 => 
                           n13871, B2 => REGISTERS_0_19_port, C1 => n13825, C2 
                           => REGISTERS_1_19_port, ZN => n15325);
   U13861 : NOR4_X1 port map( A1 => n15326, A2 => n15327, A3 => n15328, A4 => 
                           n15329, ZN => n15316);
   U13862 : OAI221_X1 port map( B1 => n11738, B2 => n365, C1 => n11002, C2 => 
                           n376, A => n15330, ZN => n15329);
   U13863 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_31_19_port, B1 => 
                           n398, B2 => REGISTERS_35_19_port, C1 => n409, C2 => 
                           REGISTERS_39_19_port, ZN => n15330);
   U13864 : OAI221_X1 port map( B1 => n11578, B2 => n420, C1 => n11706, C2 => 
                           n431, A => n15331, ZN => n15328);
   U13865 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_26_19_port, B1 => 
                           n453, B2 => REGISTERS_30_19_port, C1 => n464, C2 => 
                           REGISTERS_34_19_port, ZN => n15331);
   U13866 : OAI221_X1 port map( B1 => n11418, B2 => n475, C1 => n11546, C2 => 
                           n486, A => n15332, ZN => n15327);
   U13867 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_21_19_port, B1 => 
                           n508, B2 => REGISTERS_25_19_port, C1 => n519, C2 => 
                           REGISTERS_29_19_port, ZN => n15332);
   U13868 : OAI221_X1 port map( B1 => n11258, B2 => n530, C1 => n11386, C2 => 
                           n541, A => n15333, ZN => n15326);
   U13869 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_24_19_port, B1 => 
                           n563, B2 => REGISTERS_22_19_port, C1 => n574, C2 => 
                           REGISTERS_20_19_port, ZN => n15333);
   U13870 : AOI22_X1 port map( A1 => n13880, A2 => n5064, B1 => n13881, B2 => 
                           n5065, ZN => n15294);
   U13871 : NOR4_X1 port map( A1 => n15336, A2 => n15337, A3 => n15338, A4 => 
                           n15339, ZN => n15335);
   U13872 : OAI221_X1 port map( B1 => n11066, B2 => n310, C1 => n11002, C2 => 
                           n321, A => n15340, ZN => n15339);
   U13873 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_14_19_port, B1 => 
                           n13808, B2 => REGISTERS_38_19_port, C1 => n13889, C2
                           => REGISTERS_39_19_port, ZN => n15340);
   U13874 : OAI221_X1 port map( B1 => n10906, B2 => n13810, C1 => n10842, C2 =>
                           n13890, A => n15341, ZN => n15338);
   U13875 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_19_port, B1 => 
                           n344, B2 => REGISTERS_9_19_port, C1 => n13812, C2 =>
                           REGISTERS_16_19_port, ZN => n15341);
   U13876 : OAI221_X1 port map( B1 => n10746, B2 => n303, C1 => n10682, C2 => 
                           n13893, A => n15342, ZN => n15337);
   U13877 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_19_port, B1 => 
                           n355, B2 => REGISTERS_4_19_port, C1 => n13818, C2 =>
                           REGISTERS_11_19_port, ZN => n15342);
   U13878 : OAI221_X1 port map( B1 => n11610, B2 => n304, C1 => n10554, C2 => 
                           n13896, A => n15343, ZN => n15336);
   U13879 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_19_port, B1 => 
                           n13826, B2 => REGISTERS_0_19_port, C1 => n13824, C2 
                           => REGISTERS_6_19_port, ZN => n15343);
   U13880 : NOR4_X1 port map( A1 => n15344, A2 => n15345, A3 => n15346, A4 => 
                           n15347, ZN => n15334);
   U13881 : OAI221_X1 port map( B1 => n11674, B2 => n365, C1 => n10938, C2 => 
                           n376, A => n15348, ZN => n15347);
   U13882 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_29_19_port, B1 => 
                           n398, B2 => REGISTERS_33_19_port, C1 => n409, C2 => 
                           REGISTERS_37_19_port, ZN => n15348);
   U13883 : OAI221_X1 port map( B1 => n11514, B2 => n420, C1 => n11642, C2 => 
                           n431, A => n15349, ZN => n15346);
   U13884 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_24_19_port, B1 => 
                           n453, B2 => REGISTERS_28_19_port, C1 => n464, C2 => 
                           REGISTERS_32_19_port, ZN => n15349);
   U13885 : OAI221_X1 port map( B1 => n11354, B2 => n475, C1 => n11482, C2 => 
                           n486, A => n15350, ZN => n15345);
   U13886 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_19_19_port, B1 => 
                           n508, B2 => REGISTERS_23_19_port, C1 => n519, C2 => 
                           REGISTERS_27_19_port, ZN => n15350);
   U13887 : OAI221_X1 port map( B1 => n11194, B2 => n530, C1 => n11322, C2 => 
                           n541, A => n15351, ZN => n15344);
   U13888 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_22_19_port, B1 => 
                           n563, B2 => REGISTERS_20_19_port, C1 => n574, C2 => 
                           REGISTERS_18_19_port, ZN => n15351);
   U13889 : NOR4_X1 port map( A1 => n15354, A2 => n15355, A3 => n15356, A4 => 
                           n15357, ZN => n15353);
   U13890 : OAI221_X1 port map( B1 => n11034, B2 => n310, C1 => n10970, C2 => 
                           n321, A => n15358, ZN => n15357);
   U13891 : AOI222_X1 port map( A1 => n332, A2 => REGISTERS_13_19_port, B1 => 
                           n13808, B2 => REGISTERS_37_19_port, C1 => n13889, C2
                           => REGISTERS_38_19_port, ZN => n15358);
   U13892 : OAI221_X1 port map( B1 => n10874, B2 => n13810, C1 => n10810, C2 =>
                           n13890, A => n15359, ZN => n15356);
   U13893 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_19_port, B1 => 
                           n344, B2 => REGISTERS_8_19_port, C1 => n13812, C2 =>
                           REGISTERS_15_19_port, ZN => n15359);
   U13894 : OAI221_X1 port map( B1 => n10714, B2 => n303, C1 => n10650, C2 => 
                           n13893, A => n15360, ZN => n15355);
   U13895 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_19_port, B1 => 
                           n355, B2 => REGISTERS_3_19_port, C1 => n13818, C2 =>
                           REGISTERS_10_19_port, ZN => n15360);
   U13896 : OAI221_X1 port map( B1 => n11578, B2 => n304, C1 => n10484, C2 => 
                           n13896, A => n15361, ZN => n15354);
   U13897 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_19_port, B1 => 
                           n13917, B2 => REGISTERS_39_19_port, C1 => n13824, C2
                           => REGISTERS_5_19_port, ZN => n15361);
   U13898 : NOR4_X1 port map( A1 => n15362, A2 => n15363, A3 => n15364, A4 => 
                           n15365, ZN => n15352);
   U13899 : OAI221_X1 port map( B1 => n11642, B2 => n365, C1 => n10906, C2 => 
                           n376, A => n15366, ZN => n15365);
   U13900 : AOI222_X1 port map( A1 => n387, A2 => REGISTERS_28_19_port, B1 => 
                           n398, B2 => REGISTERS_32_19_port, C1 => n409, C2 => 
                           REGISTERS_36_19_port, ZN => n15366);
   U13901 : OAI221_X1 port map( B1 => n11482, B2 => n420, C1 => n11610, C2 => 
                           n431, A => n15367, ZN => n15364);
   U13902 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_23_19_port, B1 => 
                           n453, B2 => REGISTERS_27_19_port, C1 => n464, C2 => 
                           REGISTERS_31_19_port, ZN => n15367);
   U13903 : OAI221_X1 port map( B1 => n11322, B2 => n475, C1 => n11450, C2 => 
                           n486, A => n15368, ZN => n15363);
   U13904 : AOI222_X1 port map( A1 => n497, A2 => REGISTERS_18_19_port, B1 => 
                           n508, B2 => REGISTERS_22_19_port, C1 => n519, C2 => 
                           REGISTERS_26_19_port, ZN => n15368);
   U13905 : OAI221_X1 port map( B1 => n11162, B2 => n530, C1 => n11290, C2 => 
                           n541, A => n15369, ZN => n15362);
   U13906 : AOI222_X1 port map( A1 => n552, A2 => REGISTERS_21_19_port, B1 => 
                           n563, B2 => REGISTERS_19_19_port, C1 => n574, C2 => 
                           REGISTERS_17_19_port, ZN => n15369);
   U13907 : NAND3_X1 port map( A1 => n15370, A2 => n15371, A3 => n15372, ZN => 
                           n11884);
   U13908 : AOI221_X1 port map( B1 => n13792, B2 => n5069, C1 => n13793, C2 => 
                           MEM_IN(20), A => n15373, ZN => n15372);
   U13909 : OAI22_X1 port map( A1 => n10481, A2 => n251, B1 => n5071, B2 => 
                           n121, ZN => n15373);
   U13910 : NOR2_X1 port map( A1 => n5676, A2 => n13796, ZN => n5674);
   U13911 : INV_X1 port map( A => MEM_IN(20), ZN => n5676);
   U13912 : AOI22_X1 port map( A1 => n197, A2 => n5072, B1 => n150, B2 => n5073
                           , ZN => n15371);
   U13913 : NOR4_X1 port map( A1 => n15376, A2 => n15377, A3 => n15378, A4 => 
                           n15379, ZN => n15375);
   U13914 : OAI221_X1 port map( B1 => n11097, B2 => n309, C1 => n11033, C2 => 
                           n320, A => n15380, ZN => n15379);
   U13915 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_15_20_port, B1 => 
                           n13807, B2 => REGISTERS_11_20_port, C1 => n13808, C2
                           => REGISTERS_39_20_port, ZN => n15380);
   U13916 : OAI221_X1 port map( B1 => n10809, B2 => n13809, C1 => n10937, C2 =>
                           n13810, A => n15381, ZN => n15378);
   U13917 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_20_port, B1 =>
                           n13813, B2 => REGISTERS_6_20_port, C1 => n348, C2 =>
                           REGISTERS_10_20_port, ZN => n15381);
   U13918 : OAI221_X1 port map( B1 => n10649, B2 => n13815, C1 => n10777, C2 =>
                           n303, A => n15382, ZN => n15377);
   U13919 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_20_port, B1 =>
                           n13819, B2 => REGISTERS_2_20_port, C1 => n359, C2 =>
                           REGISTERS_5_20_port, ZN => n15382);
   U13920 : OAI221_X1 port map( B1 => n10617, B2 => n13821, C1 => n11641, C2 =>
                           n304, A => n15383, ZN => n15376);
   U13921 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_20_port, B1 => 
                           n13825, B2 => REGISTERS_0_20_port, C1 => n13826, C2 
                           => REGISTERS_1_20_port, ZN => n15383);
   U13922 : NOR4_X1 port map( A1 => n15384, A2 => n15385, A3 => n15386, A4 => 
                           n15387, ZN => n15374);
   U13923 : OAI221_X1 port map( B1 => n11705, B2 => n364, C1 => n10969, C2 => 
                           n376, A => n15388, ZN => n15387);
   U13924 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_30_20_port, B1 => 
                           n397, B2 => REGISTERS_34_20_port, C1 => n408, C2 => 
                           REGISTERS_38_20_port, ZN => n15388);
   U13925 : OAI221_X1 port map( B1 => n11545, B2 => n419, C1 => n11673, C2 => 
                           n430, A => n15389, ZN => n15386);
   U13926 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_25_20_port, B1 => 
                           n452, B2 => REGISTERS_29_20_port, C1 => n463, C2 => 
                           REGISTERS_33_20_port, ZN => n15389);
   U13927 : OAI221_X1 port map( B1 => n11385, B2 => n474, C1 => n11513, C2 => 
                           n485, A => n15390, ZN => n15385);
   U13928 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_20_20_port, B1 => 
                           n507, B2 => REGISTERS_24_20_port, C1 => n518, C2 => 
                           REGISTERS_28_20_port, ZN => n15390);
   U13929 : OAI221_X1 port map( B1 => n11225, B2 => n529, C1 => n11353, C2 => 
                           n540, A => n15391, ZN => n15384);
   U13930 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_23_20_port, B1 => 
                           n562, B2 => REGISTERS_21_20_port, C1 => n573, C2 => 
                           REGISTERS_19_20_port, ZN => n15391);
   U13931 : NOR4_X1 port map( A1 => n15394, A2 => n15395, A3 => n15396, A4 => 
                           n15397, ZN => n15393);
   U13932 : OAI221_X1 port map( B1 => n11129, B2 => n309, C1 => n11065, C2 => 
                           n320, A => n15398, ZN => n15397);
   U13933 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_16_20_port, B1 => 
                           n119, B2 => REGISTERS_14_20_port, C1 => n13807, C2 
                           => REGISTERS_12_20_port, ZN => n15398);
   U13934 : OAI221_X1 port map( B1 => n11097, B2 => n13863, C1 => n10841, C2 =>
                           n13809, A => n15399, ZN => n15396);
   U13935 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_20_port, B1 => 
                           n13865, B2 => REGISTERS_9_20_port, C1 => n13813, C2 
                           => REGISTERS_7_20_port, ZN => n15399);
   U13936 : OAI221_X1 port map( B1 => n10937, B2 => n13866, C1 => n10681, C2 =>
                           n13815, A => n15400, ZN => n15395);
   U13937 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_20_port, B1 => 
                           n13868, B2 => REGISTERS_36_20_port, C1 => n13819, C2
                           => REGISTERS_3_20_port, ZN => n15400);
   U13938 : OAI221_X1 port map( B1 => n10777, B2 => n13869, C1 => n10649, C2 =>
                           n13821, A => n15401, ZN => n15394);
   U13939 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_20_port, B1 => 
                           n13871, B2 => REGISTERS_0_20_port, C1 => n13825, C2 
                           => REGISTERS_1_20_port, ZN => n15401);
   U13940 : NOR4_X1 port map( A1 => n15402, A2 => n15403, A3 => n15404, A4 => 
                           n15405, ZN => n15392);
   U13941 : OAI221_X1 port map( B1 => n11737, B2 => n364, C1 => n11001, C2 => 
                           n375, A => n15406, ZN => n15405);
   U13942 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_31_20_port, B1 => 
                           n397, B2 => REGISTERS_35_20_port, C1 => n408, C2 => 
                           REGISTERS_39_20_port, ZN => n15406);
   U13943 : OAI221_X1 port map( B1 => n11577, B2 => n419, C1 => n11705, C2 => 
                           n430, A => n15407, ZN => n15404);
   U13944 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_26_20_port, B1 => 
                           n452, B2 => REGISTERS_30_20_port, C1 => n463, C2 => 
                           REGISTERS_34_20_port, ZN => n15407);
   U13945 : OAI221_X1 port map( B1 => n11417, B2 => n474, C1 => n11545, C2 => 
                           n485, A => n15408, ZN => n15403);
   U13946 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_21_20_port, B1 => 
                           n507, B2 => REGISTERS_25_20_port, C1 => n518, C2 => 
                           REGISTERS_29_20_port, ZN => n15408);
   U13947 : OAI221_X1 port map( B1 => n11257, B2 => n529, C1 => n11385, C2 => 
                           n540, A => n15409, ZN => n15402);
   U13948 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_24_20_port, B1 => 
                           n562, B2 => REGISTERS_22_20_port, C1 => n573, C2 => 
                           REGISTERS_20_20_port, ZN => n15409);
   U13949 : AOI22_X1 port map( A1 => n13880, A2 => n5074, B1 => n13881, B2 => 
                           n5075, ZN => n15370);
   U13950 : NOR4_X1 port map( A1 => n15412, A2 => n15413, A3 => n15414, A4 => 
                           n15415, ZN => n15411);
   U13951 : OAI221_X1 port map( B1 => n11065, B2 => n309, C1 => n11001, C2 => 
                           n320, A => n15416, ZN => n15415);
   U13952 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_14_20_port, B1 => 
                           n13808, B2 => REGISTERS_38_20_port, C1 => n13889, C2
                           => REGISTERS_39_20_port, ZN => n15416);
   U13953 : OAI221_X1 port map( B1 => n10905, B2 => n13810, C1 => n10841, C2 =>
                           n13890, A => n15417, ZN => n15414);
   U13954 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_20_port, B1 => 
                           n344, B2 => REGISTERS_9_20_port, C1 => n13812, C2 =>
                           REGISTERS_16_20_port, ZN => n15417);
   U13955 : OAI221_X1 port map( B1 => n10745, B2 => n303, C1 => n10681, C2 => 
                           n13893, A => n15418, ZN => n15413);
   U13956 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_20_port, B1 => 
                           n355, B2 => REGISTERS_4_20_port, C1 => n13818, C2 =>
                           REGISTERS_11_20_port, ZN => n15418);
   U13957 : OAI221_X1 port map( B1 => n11609, B2 => n304, C1 => n10553, C2 => 
                           n13896, A => n15419, ZN => n15412);
   U13958 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_20_port, B1 => 
                           n13826, B2 => REGISTERS_0_20_port, C1 => n13824, C2 
                           => REGISTERS_6_20_port, ZN => n15419);
   U13959 : NOR4_X1 port map( A1 => n15420, A2 => n15421, A3 => n15422, A4 => 
                           n15423, ZN => n15410);
   U13960 : OAI221_X1 port map( B1 => n11673, B2 => n364, C1 => n10937, C2 => 
                           n375, A => n15424, ZN => n15423);
   U13961 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_29_20_port, B1 => 
                           n397, B2 => REGISTERS_33_20_port, C1 => n408, C2 => 
                           REGISTERS_37_20_port, ZN => n15424);
   U13962 : OAI221_X1 port map( B1 => n11513, B2 => n419, C1 => n11641, C2 => 
                           n430, A => n15425, ZN => n15422);
   U13963 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_24_20_port, B1 => 
                           n452, B2 => REGISTERS_28_20_port, C1 => n463, C2 => 
                           REGISTERS_32_20_port, ZN => n15425);
   U13964 : OAI221_X1 port map( B1 => n11353, B2 => n474, C1 => n11481, C2 => 
                           n485, A => n15426, ZN => n15421);
   U13965 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_19_20_port, B1 => 
                           n507, B2 => REGISTERS_23_20_port, C1 => n518, C2 => 
                           REGISTERS_27_20_port, ZN => n15426);
   U13966 : OAI221_X1 port map( B1 => n11193, B2 => n529, C1 => n11321, C2 => 
                           n540, A => n15427, ZN => n15420);
   U13967 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_22_20_port, B1 => 
                           n562, B2 => REGISTERS_20_20_port, C1 => n573, C2 => 
                           REGISTERS_18_20_port, ZN => n15427);
   U13968 : NOR4_X1 port map( A1 => n15430, A2 => n15431, A3 => n15432, A4 => 
                           n15433, ZN => n15429);
   U13969 : OAI221_X1 port map( B1 => n11033, B2 => n309, C1 => n10969, C2 => 
                           n320, A => n15434, ZN => n15433);
   U13970 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_13_20_port, B1 => 
                           n13808, B2 => REGISTERS_37_20_port, C1 => n13889, C2
                           => REGISTERS_38_20_port, ZN => n15434);
   U13971 : OAI221_X1 port map( B1 => n10873, B2 => n13810, C1 => n10809, C2 =>
                           n13890, A => n15435, ZN => n15432);
   U13972 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_20_port, B1 => 
                           n344, B2 => REGISTERS_8_20_port, C1 => n13812, C2 =>
                           REGISTERS_15_20_port, ZN => n15435);
   U13973 : OAI221_X1 port map( B1 => n10713, B2 => n303, C1 => n10649, C2 => 
                           n13893, A => n15436, ZN => n15431);
   U13974 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_20_port, B1 => 
                           n355, B2 => REGISTERS_3_20_port, C1 => n13818, C2 =>
                           REGISTERS_10_20_port, ZN => n15436);
   U13975 : OAI221_X1 port map( B1 => n11577, B2 => n304, C1 => n10481, C2 => 
                           n13896, A => n15437, ZN => n15430);
   U13976 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_20_port, B1 => 
                           n13917, B2 => REGISTERS_39_20_port, C1 => n13824, C2
                           => REGISTERS_5_20_port, ZN => n15437);
   U13977 : NOR4_X1 port map( A1 => n15438, A2 => n15439, A3 => n15440, A4 => 
                           n15441, ZN => n15428);
   U13978 : OAI221_X1 port map( B1 => n11641, B2 => n364, C1 => n10905, C2 => 
                           n375, A => n15442, ZN => n15441);
   U13979 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_28_20_port, B1 => 
                           n397, B2 => REGISTERS_32_20_port, C1 => n408, C2 => 
                           REGISTERS_36_20_port, ZN => n15442);
   U13980 : OAI221_X1 port map( B1 => n11481, B2 => n419, C1 => n11609, C2 => 
                           n430, A => n15443, ZN => n15440);
   U13981 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_23_20_port, B1 => 
                           n452, B2 => REGISTERS_27_20_port, C1 => n463, C2 => 
                           REGISTERS_31_20_port, ZN => n15443);
   U13982 : OAI221_X1 port map( B1 => n11321, B2 => n474, C1 => n11449, C2 => 
                           n485, A => n15444, ZN => n15439);
   U13983 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_18_20_port, B1 => 
                           n507, B2 => REGISTERS_22_20_port, C1 => n518, C2 => 
                           REGISTERS_26_20_port, ZN => n15444);
   U13984 : OAI221_X1 port map( B1 => n11161, B2 => n529, C1 => n11289, C2 => 
                           n540, A => n15445, ZN => n15438);
   U13985 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_21_20_port, B1 => 
                           n562, B2 => REGISTERS_19_20_port, C1 => n573, C2 => 
                           REGISTERS_17_20_port, ZN => n15445);
   U13986 : NAND3_X1 port map( A1 => n15446, A2 => n15447, A3 => n15448, ZN => 
                           n11883);
   U13987 : AOI221_X1 port map( B1 => n13792, B2 => n5079, C1 => n13793, C2 => 
                           MEM_IN(21), A => n15449, ZN => n15448);
   U13988 : OAI22_X1 port map( A1 => n10478, A2 => n251, B1 => n5081, B2 => 
                           n121, ZN => n15449);
   U13989 : NOR2_X1 port map( A1 => n5683, A2 => n13796, ZN => n5681);
   U13990 : INV_X1 port map( A => MEM_IN(21), ZN => n5683);
   U13991 : AOI22_X1 port map( A1 => n197, A2 => n5082, B1 => n150, B2 => n5083
                           , ZN => n15447);
   U13992 : NOR4_X1 port map( A1 => n15452, A2 => n15453, A3 => n15454, A4 => 
                           n15455, ZN => n15451);
   U13993 : OAI221_X1 port map( B1 => n11096, B2 => n309, C1 => n11032, C2 => 
                           n320, A => n15456, ZN => n15455);
   U13994 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_15_21_port, B1 => 
                           n13807, B2 => REGISTERS_11_21_port, C1 => n13808, C2
                           => REGISTERS_39_21_port, ZN => n15456);
   U13995 : OAI221_X1 port map( B1 => n10808, B2 => n13809, C1 => n10936, C2 =>
                           n13810, A => n15457, ZN => n15454);
   U13996 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_21_port, B1 =>
                           n13813, B2 => REGISTERS_6_21_port, C1 => n348, C2 =>
                           REGISTERS_10_21_port, ZN => n15457);
   U13997 : OAI221_X1 port map( B1 => n10648, B2 => n13815, C1 => n10776, C2 =>
                           n303, A => n15458, ZN => n15453);
   U13998 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_21_port, B1 =>
                           n13819, B2 => REGISTERS_2_21_port, C1 => n359, C2 =>
                           REGISTERS_5_21_port, ZN => n15458);
   U13999 : OAI221_X1 port map( B1 => n10616, B2 => n13821, C1 => n11640, C2 =>
                           n304, A => n15459, ZN => n15452);
   U14000 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_21_port, B1 => 
                           n13825, B2 => REGISTERS_0_21_port, C1 => n13826, C2 
                           => REGISTERS_1_21_port, ZN => n15459);
   U14001 : NOR4_X1 port map( A1 => n15460, A2 => n15461, A3 => n15462, A4 => 
                           n15463, ZN => n15450);
   U14002 : OAI221_X1 port map( B1 => n11704, B2 => n364, C1 => n10968, C2 => 
                           n375, A => n15464, ZN => n15463);
   U14003 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_30_21_port, B1 => 
                           n397, B2 => REGISTERS_34_21_port, C1 => n408, C2 => 
                           REGISTERS_38_21_port, ZN => n15464);
   U14004 : OAI221_X1 port map( B1 => n11544, B2 => n419, C1 => n11672, C2 => 
                           n430, A => n15465, ZN => n15462);
   U14005 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_25_21_port, B1 => 
                           n452, B2 => REGISTERS_29_21_port, C1 => n463, C2 => 
                           REGISTERS_33_21_port, ZN => n15465);
   U14006 : OAI221_X1 port map( B1 => n11384, B2 => n474, C1 => n11512, C2 => 
                           n485, A => n15466, ZN => n15461);
   U14007 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_20_21_port, B1 => 
                           n507, B2 => REGISTERS_24_21_port, C1 => n518, C2 => 
                           REGISTERS_28_21_port, ZN => n15466);
   U14008 : OAI221_X1 port map( B1 => n11224, B2 => n529, C1 => n11352, C2 => 
                           n540, A => n15467, ZN => n15460);
   U14009 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_23_21_port, B1 => 
                           n562, B2 => REGISTERS_21_21_port, C1 => n573, C2 => 
                           REGISTERS_19_21_port, ZN => n15467);
   U14010 : NOR4_X1 port map( A1 => n15470, A2 => n15471, A3 => n15472, A4 => 
                           n15473, ZN => n15469);
   U14011 : OAI221_X1 port map( B1 => n11128, B2 => n309, C1 => n11064, C2 => 
                           n320, A => n15474, ZN => n15473);
   U14012 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_16_21_port, B1 => 
                           n119, B2 => REGISTERS_14_21_port, C1 => n13807, C2 
                           => REGISTERS_12_21_port, ZN => n15474);
   U14013 : OAI221_X1 port map( B1 => n11096, B2 => n13863, C1 => n10840, C2 =>
                           n13809, A => n15475, ZN => n15472);
   U14014 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_21_port, B1 => 
                           n13865, B2 => REGISTERS_9_21_port, C1 => n13813, C2 
                           => REGISTERS_7_21_port, ZN => n15475);
   U14015 : OAI221_X1 port map( B1 => n10936, B2 => n13866, C1 => n10680, C2 =>
                           n13815, A => n15476, ZN => n15471);
   U14016 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_21_port, B1 => 
                           n13868, B2 => REGISTERS_36_21_port, C1 => n13819, C2
                           => REGISTERS_3_21_port, ZN => n15476);
   U14017 : OAI221_X1 port map( B1 => n10776, B2 => n13869, C1 => n10648, C2 =>
                           n13821, A => n15477, ZN => n15470);
   U14018 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_21_port, B1 => 
                           n13871, B2 => REGISTERS_0_21_port, C1 => n13825, C2 
                           => REGISTERS_1_21_port, ZN => n15477);
   U14019 : NOR4_X1 port map( A1 => n15478, A2 => n15479, A3 => n15480, A4 => 
                           n15481, ZN => n15468);
   U14020 : OAI221_X1 port map( B1 => n11736, B2 => n364, C1 => n11000, C2 => 
                           n375, A => n15482, ZN => n15481);
   U14021 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_31_21_port, B1 => 
                           n397, B2 => REGISTERS_35_21_port, C1 => n408, C2 => 
                           REGISTERS_39_21_port, ZN => n15482);
   U14022 : OAI221_X1 port map( B1 => n11576, B2 => n419, C1 => n11704, C2 => 
                           n430, A => n15483, ZN => n15480);
   U14023 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_26_21_port, B1 => 
                           n452, B2 => REGISTERS_30_21_port, C1 => n463, C2 => 
                           REGISTERS_34_21_port, ZN => n15483);
   U14024 : OAI221_X1 port map( B1 => n11416, B2 => n474, C1 => n11544, C2 => 
                           n485, A => n15484, ZN => n15479);
   U14025 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_21_21_port, B1 => 
                           n507, B2 => REGISTERS_25_21_port, C1 => n518, C2 => 
                           REGISTERS_29_21_port, ZN => n15484);
   U14026 : OAI221_X1 port map( B1 => n11256, B2 => n529, C1 => n11384, C2 => 
                           n540, A => n15485, ZN => n15478);
   U14027 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_24_21_port, B1 => 
                           n562, B2 => REGISTERS_22_21_port, C1 => n573, C2 => 
                           REGISTERS_20_21_port, ZN => n15485);
   U14028 : AOI22_X1 port map( A1 => n13880, A2 => n5084, B1 => n13881, B2 => 
                           n5085, ZN => n15446);
   U14029 : NOR4_X1 port map( A1 => n15488, A2 => n15489, A3 => n15490, A4 => 
                           n15491, ZN => n15487);
   U14030 : OAI221_X1 port map( B1 => n11064, B2 => n309, C1 => n11000, C2 => 
                           n320, A => n15492, ZN => n15491);
   U14031 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_14_21_port, B1 => 
                           n13808, B2 => REGISTERS_38_21_port, C1 => n13889, C2
                           => REGISTERS_39_21_port, ZN => n15492);
   U14032 : OAI221_X1 port map( B1 => n10904, B2 => n13810, C1 => n10840, C2 =>
                           n13890, A => n15493, ZN => n15490);
   U14033 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_21_port, B1 => 
                           n345, B2 => REGISTERS_9_21_port, C1 => n13812, C2 =>
                           REGISTERS_16_21_port, ZN => n15493);
   U14034 : OAI221_X1 port map( B1 => n10744, B2 => n303, C1 => n10680, C2 => 
                           n13893, A => n15494, ZN => n15489);
   U14035 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_21_port, B1 => 
                           n356, B2 => REGISTERS_4_21_port, C1 => n13818, C2 =>
                           REGISTERS_11_21_port, ZN => n15494);
   U14036 : OAI221_X1 port map( B1 => n11608, B2 => n304, C1 => n10552, C2 => 
                           n13896, A => n15495, ZN => n15488);
   U14037 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_21_port, B1 => 
                           n13826, B2 => REGISTERS_0_21_port, C1 => n13824, C2 
                           => REGISTERS_6_21_port, ZN => n15495);
   U14038 : NOR4_X1 port map( A1 => n15496, A2 => n15497, A3 => n15498, A4 => 
                           n15499, ZN => n15486);
   U14039 : OAI221_X1 port map( B1 => n11672, B2 => n364, C1 => n10936, C2 => 
                           n375, A => n15500, ZN => n15499);
   U14040 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_29_21_port, B1 => 
                           n397, B2 => REGISTERS_33_21_port, C1 => n408, C2 => 
                           REGISTERS_37_21_port, ZN => n15500);
   U14041 : OAI221_X1 port map( B1 => n11512, B2 => n419, C1 => n11640, C2 => 
                           n430, A => n15501, ZN => n15498);
   U14042 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_24_21_port, B1 => 
                           n452, B2 => REGISTERS_28_21_port, C1 => n463, C2 => 
                           REGISTERS_32_21_port, ZN => n15501);
   U14043 : OAI221_X1 port map( B1 => n11352, B2 => n474, C1 => n11480, C2 => 
                           n485, A => n15502, ZN => n15497);
   U14044 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_19_21_port, B1 => 
                           n507, B2 => REGISTERS_23_21_port, C1 => n518, C2 => 
                           REGISTERS_27_21_port, ZN => n15502);
   U14045 : OAI221_X1 port map( B1 => n11192, B2 => n529, C1 => n11320, C2 => 
                           n540, A => n15503, ZN => n15496);
   U14046 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_22_21_port, B1 => 
                           n562, B2 => REGISTERS_20_21_port, C1 => n573, C2 => 
                           REGISTERS_18_21_port, ZN => n15503);
   U14047 : NOR4_X1 port map( A1 => n15506, A2 => n15507, A3 => n15508, A4 => 
                           n15509, ZN => n15505);
   U14048 : OAI221_X1 port map( B1 => n11032, B2 => n309, C1 => n10968, C2 => 
                           n320, A => n15510, ZN => n15509);
   U14049 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_13_21_port, B1 => 
                           n13808, B2 => REGISTERS_37_21_port, C1 => n13889, C2
                           => REGISTERS_38_21_port, ZN => n15510);
   U14050 : OAI221_X1 port map( B1 => n10872, B2 => n13810, C1 => n10808, C2 =>
                           n13890, A => n15511, ZN => n15508);
   U14051 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_21_port, B1 => 
                           n344, B2 => REGISTERS_8_21_port, C1 => n13812, C2 =>
                           REGISTERS_15_21_port, ZN => n15511);
   U14052 : OAI221_X1 port map( B1 => n10712, B2 => n303, C1 => n10648, C2 => 
                           n13893, A => n15512, ZN => n15507);
   U14053 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_21_port, B1 => 
                           n355, B2 => REGISTERS_3_21_port, C1 => n13818, C2 =>
                           REGISTERS_10_21_port, ZN => n15512);
   U14054 : OAI221_X1 port map( B1 => n11576, B2 => n304, C1 => n10478, C2 => 
                           n13896, A => n15513, ZN => n15506);
   U14055 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_21_port, B1 => 
                           n13917, B2 => REGISTERS_39_21_port, C1 => n13824, C2
                           => REGISTERS_5_21_port, ZN => n15513);
   U14056 : NOR4_X1 port map( A1 => n15514, A2 => n15515, A3 => n15516, A4 => 
                           n15517, ZN => n15504);
   U14057 : OAI221_X1 port map( B1 => n11640, B2 => n364, C1 => n10904, C2 => 
                           n375, A => n15518, ZN => n15517);
   U14058 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_28_21_port, B1 => 
                           n397, B2 => REGISTERS_32_21_port, C1 => n408, C2 => 
                           REGISTERS_36_21_port, ZN => n15518);
   U14059 : OAI221_X1 port map( B1 => n11480, B2 => n419, C1 => n11608, C2 => 
                           n430, A => n15519, ZN => n15516);
   U14060 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_23_21_port, B1 => 
                           n452, B2 => REGISTERS_27_21_port, C1 => n463, C2 => 
                           REGISTERS_31_21_port, ZN => n15519);
   U14061 : OAI221_X1 port map( B1 => n11320, B2 => n474, C1 => n11448, C2 => 
                           n485, A => n15520, ZN => n15515);
   U14062 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_18_21_port, B1 => 
                           n507, B2 => REGISTERS_22_21_port, C1 => n518, C2 => 
                           REGISTERS_26_21_port, ZN => n15520);
   U14063 : OAI221_X1 port map( B1 => n11160, B2 => n529, C1 => n11288, C2 => 
                           n540, A => n15521, ZN => n15514);
   U14064 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_21_21_port, B1 => 
                           n562, B2 => REGISTERS_19_21_port, C1 => n573, C2 => 
                           REGISTERS_17_21_port, ZN => n15521);
   U14065 : NAND3_X1 port map( A1 => n15522, A2 => n15523, A3 => n15524, ZN => 
                           n11882);
   U14066 : AOI221_X1 port map( B1 => n13792, B2 => n5089, C1 => n13793, C2 => 
                           MEM_IN(22), A => n15525, ZN => n15524);
   U14067 : OAI22_X1 port map( A1 => n10475, A2 => n251, B1 => n5091, B2 => 
                           n121, ZN => n15525);
   U14068 : NOR2_X1 port map( A1 => n5690, A2 => n13796, ZN => n5688);
   U14069 : INV_X1 port map( A => MEM_IN(22), ZN => n5690);
   U14070 : AOI22_X1 port map( A1 => n197, A2 => n5092, B1 => n150, B2 => n5093
                           , ZN => n15523);
   U14071 : NOR4_X1 port map( A1 => n15528, A2 => n15529, A3 => n15530, A4 => 
                           n15531, ZN => n15527);
   U14072 : OAI221_X1 port map( B1 => n11095, B2 => n309, C1 => n11031, C2 => 
                           n320, A => n15532, ZN => n15531);
   U14073 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_15_22_port, B1 => 
                           n13807, B2 => REGISTERS_11_22_port, C1 => n13808, C2
                           => REGISTERS_39_22_port, ZN => n15532);
   U14074 : OAI221_X1 port map( B1 => n10807, B2 => n13809, C1 => n10935, C2 =>
                           n13810, A => n15533, ZN => n15530);
   U14075 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_22_port, B1 =>
                           n13813, B2 => REGISTERS_6_22_port, C1 => n348, C2 =>
                           REGISTERS_10_22_port, ZN => n15533);
   U14076 : OAI221_X1 port map( B1 => n10647, B2 => n13815, C1 => n10775, C2 =>
                           n303, A => n15534, ZN => n15529);
   U14077 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_22_port, B1 =>
                           n13819, B2 => REGISTERS_2_22_port, C1 => n359, C2 =>
                           REGISTERS_5_22_port, ZN => n15534);
   U14078 : OAI221_X1 port map( B1 => n10615, B2 => n13821, C1 => n11639, C2 =>
                           n304, A => n15535, ZN => n15528);
   U14079 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_22_port, B1 => 
                           n13825, B2 => REGISTERS_0_22_port, C1 => n13826, C2 
                           => REGISTERS_1_22_port, ZN => n15535);
   U14080 : NOR4_X1 port map( A1 => n15536, A2 => n15537, A3 => n15538, A4 => 
                           n15539, ZN => n15526);
   U14081 : OAI221_X1 port map( B1 => n11703, B2 => n364, C1 => n10967, C2 => 
                           n375, A => n15540, ZN => n15539);
   U14082 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_30_22_port, B1 => 
                           n397, B2 => REGISTERS_34_22_port, C1 => n408, C2 => 
                           REGISTERS_38_22_port, ZN => n15540);
   U14083 : OAI221_X1 port map( B1 => n11543, B2 => n419, C1 => n11671, C2 => 
                           n430, A => n15541, ZN => n15538);
   U14084 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_25_22_port, B1 => 
                           n452, B2 => REGISTERS_29_22_port, C1 => n463, C2 => 
                           REGISTERS_33_22_port, ZN => n15541);
   U14085 : OAI221_X1 port map( B1 => n11383, B2 => n474, C1 => n11511, C2 => 
                           n485, A => n15542, ZN => n15537);
   U14086 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_20_22_port, B1 => 
                           n507, B2 => REGISTERS_24_22_port, C1 => n518, C2 => 
                           REGISTERS_28_22_port, ZN => n15542);
   U14087 : OAI221_X1 port map( B1 => n11223, B2 => n529, C1 => n11351, C2 => 
                           n540, A => n15543, ZN => n15536);
   U14088 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_23_22_port, B1 => 
                           n562, B2 => REGISTERS_21_22_port, C1 => n573, C2 => 
                           REGISTERS_19_22_port, ZN => n15543);
   U14089 : NOR4_X1 port map( A1 => n15546, A2 => n15547, A3 => n15548, A4 => 
                           n15549, ZN => n15545);
   U14090 : OAI221_X1 port map( B1 => n11127, B2 => n309, C1 => n11063, C2 => 
                           n320, A => n15550, ZN => n15549);
   U14091 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_16_22_port, B1 => 
                           n119, B2 => REGISTERS_14_22_port, C1 => n13807, C2 
                           => REGISTERS_12_22_port, ZN => n15550);
   U14092 : OAI221_X1 port map( B1 => n11095, B2 => n13863, C1 => n10839, C2 =>
                           n13809, A => n15551, ZN => n15548);
   U14093 : AOI222_X1 port map( A1 => n341, A2 => REGISTERS_11_22_port, B1 => 
                           n13865, B2 => REGISTERS_9_22_port, C1 => n13813, C2 
                           => REGISTERS_7_22_port, ZN => n15551);
   U14094 : OAI221_X1 port map( B1 => n10935, B2 => n13866, C1 => n10679, C2 =>
                           n13815, A => n15552, ZN => n15547);
   U14095 : AOI222_X1 port map( A1 => n352, A2 => REGISTERS_6_22_port, B1 => 
                           n13868, B2 => REGISTERS_36_22_port, C1 => n13819, C2
                           => REGISTERS_3_22_port, ZN => n15552);
   U14096 : OAI221_X1 port map( B1 => n10775, B2 => n13869, C1 => n10647, C2 =>
                           n13821, A => n15553, ZN => n15546);
   U14097 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_22_port, B1 => 
                           n13871, B2 => REGISTERS_0_22_port, C1 => n13825, C2 
                           => REGISTERS_1_22_port, ZN => n15553);
   U14098 : NOR4_X1 port map( A1 => n15554, A2 => n15555, A3 => n15556, A4 => 
                           n15557, ZN => n15544);
   U14099 : OAI221_X1 port map( B1 => n11735, B2 => n364, C1 => n10999, C2 => 
                           n375, A => n15558, ZN => n15557);
   U14100 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_31_22_port, B1 => 
                           n397, B2 => REGISTERS_35_22_port, C1 => n408, C2 => 
                           REGISTERS_39_22_port, ZN => n15558);
   U14101 : OAI221_X1 port map( B1 => n11575, B2 => n419, C1 => n11703, C2 => 
                           n430, A => n15559, ZN => n15556);
   U14102 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_26_22_port, B1 => 
                           n452, B2 => REGISTERS_30_22_port, C1 => n463, C2 => 
                           REGISTERS_34_22_port, ZN => n15559);
   U14103 : OAI221_X1 port map( B1 => n11415, B2 => n474, C1 => n11543, C2 => 
                           n485, A => n15560, ZN => n15555);
   U14104 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_21_22_port, B1 => 
                           n507, B2 => REGISTERS_25_22_port, C1 => n518, C2 => 
                           REGISTERS_29_22_port, ZN => n15560);
   U14105 : OAI221_X1 port map( B1 => n11255, B2 => n529, C1 => n11383, C2 => 
                           n540, A => n15561, ZN => n15554);
   U14106 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_24_22_port, B1 => 
                           n562, B2 => REGISTERS_22_22_port, C1 => n573, C2 => 
                           REGISTERS_20_22_port, ZN => n15561);
   U14107 : AOI22_X1 port map( A1 => n13880, A2 => n5094, B1 => n13881, B2 => 
                           n5095, ZN => n15522);
   U14108 : NOR4_X1 port map( A1 => n15564, A2 => n15565, A3 => n15566, A4 => 
                           n15567, ZN => n15563);
   U14109 : OAI221_X1 port map( B1 => n11063, B2 => n309, C1 => n10999, C2 => 
                           n320, A => n15568, ZN => n15567);
   U14110 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_14_22_port, B1 => 
                           n13808, B2 => REGISTERS_38_22_port, C1 => n13889, C2
                           => REGISTERS_39_22_port, ZN => n15568);
   U14111 : OAI221_X1 port map( B1 => n10903, B2 => n13810, C1 => n10839, C2 =>
                           n13890, A => n15569, ZN => n15566);
   U14112 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_22_port, B1 => 
                           n345, B2 => REGISTERS_9_22_port, C1 => n13812, C2 =>
                           REGISTERS_16_22_port, ZN => n15569);
   U14113 : OAI221_X1 port map( B1 => n10743, B2 => n303, C1 => n10679, C2 => 
                           n13893, A => n15570, ZN => n15565);
   U14114 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_22_port, B1 => 
                           n356, B2 => REGISTERS_4_22_port, C1 => n13818, C2 =>
                           REGISTERS_11_22_port, ZN => n15570);
   U14115 : OAI221_X1 port map( B1 => n11607, B2 => n304, C1 => n10551, C2 => 
                           n13896, A => n15571, ZN => n15564);
   U14116 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_22_port, B1 => 
                           n13826, B2 => REGISTERS_0_22_port, C1 => n13824, C2 
                           => REGISTERS_6_22_port, ZN => n15571);
   U14117 : NOR4_X1 port map( A1 => n15572, A2 => n15573, A3 => n15574, A4 => 
                           n15575, ZN => n15562);
   U14118 : OAI221_X1 port map( B1 => n11671, B2 => n364, C1 => n10935, C2 => 
                           n375, A => n15576, ZN => n15575);
   U14119 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_29_22_port, B1 => 
                           n397, B2 => REGISTERS_33_22_port, C1 => n408, C2 => 
                           REGISTERS_37_22_port, ZN => n15576);
   U14120 : OAI221_X1 port map( B1 => n11511, B2 => n419, C1 => n11639, C2 => 
                           n430, A => n15577, ZN => n15574);
   U14121 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_24_22_port, B1 => 
                           n452, B2 => REGISTERS_28_22_port, C1 => n463, C2 => 
                           REGISTERS_32_22_port, ZN => n15577);
   U14122 : OAI221_X1 port map( B1 => n11351, B2 => n474, C1 => n11479, C2 => 
                           n485, A => n15578, ZN => n15573);
   U14123 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_19_22_port, B1 => 
                           n507, B2 => REGISTERS_23_22_port, C1 => n518, C2 => 
                           REGISTERS_27_22_port, ZN => n15578);
   U14124 : OAI221_X1 port map( B1 => n11191, B2 => n529, C1 => n11319, C2 => 
                           n540, A => n15579, ZN => n15572);
   U14125 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_22_22_port, B1 => 
                           n562, B2 => REGISTERS_20_22_port, C1 => n573, C2 => 
                           REGISTERS_18_22_port, ZN => n15579);
   U14126 : NOR4_X1 port map( A1 => n15582, A2 => n15583, A3 => n15584, A4 => 
                           n15585, ZN => n15581);
   U14127 : OAI221_X1 port map( B1 => n11031, B2 => n309, C1 => n10967, C2 => 
                           n320, A => n15586, ZN => n15585);
   U14128 : AOI222_X1 port map( A1 => n331, A2 => REGISTERS_13_22_port, B1 => 
                           n13808, B2 => REGISTERS_37_22_port, C1 => n13889, C2
                           => REGISTERS_38_22_port, ZN => n15586);
   U14129 : OAI221_X1 port map( B1 => n10871, B2 => n13810, C1 => n10807, C2 =>
                           n13890, A => n15587, ZN => n15584);
   U14130 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_22_port, B1 => 
                           n345, B2 => REGISTERS_8_22_port, C1 => n13812, C2 =>
                           REGISTERS_15_22_port, ZN => n15587);
   U14131 : OAI221_X1 port map( B1 => n10711, B2 => n303, C1 => n10647, C2 => 
                           n13893, A => n15588, ZN => n15583);
   U14132 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_22_port, B1 => 
                           n356, B2 => REGISTERS_3_22_port, C1 => n13818, C2 =>
                           REGISTERS_10_22_port, ZN => n15588);
   U14133 : OAI221_X1 port map( B1 => n11575, B2 => n304, C1 => n10475, C2 => 
                           n13896, A => n15589, ZN => n15582);
   U14134 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_22_port, B1 => 
                           n13917, B2 => REGISTERS_39_22_port, C1 => n13824, C2
                           => REGISTERS_5_22_port, ZN => n15589);
   U14135 : NOR4_X1 port map( A1 => n15590, A2 => n15591, A3 => n15592, A4 => 
                           n15593, ZN => n15580);
   U14136 : OAI221_X1 port map( B1 => n11639, B2 => n364, C1 => n10903, C2 => 
                           n375, A => n15594, ZN => n15593);
   U14137 : AOI222_X1 port map( A1 => n386, A2 => REGISTERS_28_22_port, B1 => 
                           n397, B2 => REGISTERS_32_22_port, C1 => n408, C2 => 
                           REGISTERS_36_22_port, ZN => n15594);
   U14138 : OAI221_X1 port map( B1 => n11479, B2 => n419, C1 => n11607, C2 => 
                           n430, A => n15595, ZN => n15592);
   U14139 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_23_22_port, B1 => 
                           n452, B2 => REGISTERS_27_22_port, C1 => n463, C2 => 
                           REGISTERS_31_22_port, ZN => n15595);
   U14140 : OAI221_X1 port map( B1 => n11319, B2 => n474, C1 => n11447, C2 => 
                           n485, A => n15596, ZN => n15591);
   U14141 : AOI222_X1 port map( A1 => n496, A2 => REGISTERS_18_22_port, B1 => 
                           n507, B2 => REGISTERS_22_22_port, C1 => n518, C2 => 
                           REGISTERS_26_22_port, ZN => n15596);
   U14142 : OAI221_X1 port map( B1 => n11159, B2 => n529, C1 => n11287, C2 => 
                           n540, A => n15597, ZN => n15590);
   U14143 : AOI222_X1 port map( A1 => n551, A2 => REGISTERS_21_22_port, B1 => 
                           n562, B2 => REGISTERS_19_22_port, C1 => n573, C2 => 
                           REGISTERS_17_22_port, ZN => n15597);
   U14144 : NAND3_X1 port map( A1 => n15598, A2 => n15599, A3 => n15600, ZN => 
                           n11881);
   U14145 : AOI221_X1 port map( B1 => n13792, B2 => n5099, C1 => n13793, C2 => 
                           MEM_IN(23), A => n15601, ZN => n15600);
   U14146 : OAI22_X1 port map( A1 => n10472, A2 => n251, B1 => n5101, B2 => 
                           n121, ZN => n15601);
   U14147 : NOR2_X1 port map( A1 => n5697, A2 => n13796, ZN => n5695);
   U14148 : INV_X1 port map( A => MEM_IN(23), ZN => n5697);
   U14149 : AOI22_X1 port map( A1 => n197, A2 => n5102, B1 => n150, B2 => n5103
                           , ZN => n15599);
   U14150 : NOR4_X1 port map( A1 => n15604, A2 => n15605, A3 => n15606, A4 => 
                           n15607, ZN => n15603);
   U14151 : OAI221_X1 port map( B1 => n11094, B2 => n308, C1 => n11030, C2 => 
                           n319, A => n15608, ZN => n15607);
   U14152 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_15_23_port, B1 => 
                           n13807, B2 => REGISTERS_11_23_port, C1 => n13808, C2
                           => REGISTERS_39_23_port, ZN => n15608);
   U14153 : OAI221_X1 port map( B1 => n10806, B2 => n13809, C1 => n10934, C2 =>
                           n13810, A => n15609, ZN => n15606);
   U14154 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_23_port, B1 =>
                           n13813, B2 => REGISTERS_6_23_port, C1 => n349, C2 =>
                           REGISTERS_10_23_port, ZN => n15609);
   U14155 : OAI221_X1 port map( B1 => n10646, B2 => n13815, C1 => n10774, C2 =>
                           n303, A => n15610, ZN => n15605);
   U14156 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_23_port, B1 =>
                           n13819, B2 => REGISTERS_2_23_port, C1 => n360, C2 =>
                           REGISTERS_5_23_port, ZN => n15610);
   U14157 : OAI221_X1 port map( B1 => n10614, B2 => n13821, C1 => n11638, C2 =>
                           n304, A => n15611, ZN => n15604);
   U14158 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_23_port, B1 => 
                           n13825, B2 => REGISTERS_0_23_port, C1 => n13826, C2 
                           => REGISTERS_1_23_port, ZN => n15611);
   U14159 : NOR4_X1 port map( A1 => n15612, A2 => n15613, A3 => n15614, A4 => 
                           n15615, ZN => n15602);
   U14160 : OAI221_X1 port map( B1 => n11702, B2 => n363, C1 => n10966, C2 => 
                           n375, A => n15616, ZN => n15615);
   U14161 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_30_23_port, B1 => 
                           n396, B2 => REGISTERS_34_23_port, C1 => n407, C2 => 
                           REGISTERS_38_23_port, ZN => n15616);
   U14162 : OAI221_X1 port map( B1 => n11542, B2 => n418, C1 => n11670, C2 => 
                           n429, A => n15617, ZN => n15614);
   U14163 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_25_23_port, B1 => 
                           n451, B2 => REGISTERS_29_23_port, C1 => n462, C2 => 
                           REGISTERS_33_23_port, ZN => n15617);
   U14164 : OAI221_X1 port map( B1 => n11382, B2 => n473, C1 => n11510, C2 => 
                           n484, A => n15618, ZN => n15613);
   U14165 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_20_23_port, B1 => 
                           n506, B2 => REGISTERS_24_23_port, C1 => n517, C2 => 
                           REGISTERS_28_23_port, ZN => n15618);
   U14166 : OAI221_X1 port map( B1 => n11222, B2 => n528, C1 => n11350, C2 => 
                           n539, A => n15619, ZN => n15612);
   U14167 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_23_23_port, B1 => 
                           n561, B2 => REGISTERS_21_23_port, C1 => n572, C2 => 
                           REGISTERS_19_23_port, ZN => n15619);
   U14168 : NOR4_X1 port map( A1 => n15622, A2 => n15623, A3 => n15624, A4 => 
                           n15625, ZN => n15621);
   U14169 : OAI221_X1 port map( B1 => n11126, B2 => n308, C1 => n11062, C2 => 
                           n319, A => n15626, ZN => n15625);
   U14170 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_16_23_port, B1 => 
                           n119, B2 => REGISTERS_14_23_port, C1 => n13807, C2 
                           => REGISTERS_12_23_port, ZN => n15626);
   U14171 : OAI221_X1 port map( B1 => n11094, B2 => n13863, C1 => n10838, C2 =>
                           n13809, A => n15627, ZN => n15624);
   U14172 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_23_port, B1 => 
                           n13865, B2 => REGISTERS_9_23_port, C1 => n13813, C2 
                           => REGISTERS_7_23_port, ZN => n15627);
   U14173 : OAI221_X1 port map( B1 => n10934, B2 => n13866, C1 => n10678, C2 =>
                           n13815, A => n15628, ZN => n15623);
   U14174 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_23_port, B1 => 
                           n13868, B2 => REGISTERS_36_23_port, C1 => n13819, C2
                           => REGISTERS_3_23_port, ZN => n15628);
   U14175 : OAI221_X1 port map( B1 => n10774, B2 => n13869, C1 => n10646, C2 =>
                           n13821, A => n15629, ZN => n15622);
   U14176 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_23_port, B1 => 
                           n13871, B2 => REGISTERS_0_23_port, C1 => n13825, C2 
                           => REGISTERS_1_23_port, ZN => n15629);
   U14177 : NOR4_X1 port map( A1 => n15630, A2 => n15631, A3 => n15632, A4 => 
                           n15633, ZN => n15620);
   U14178 : OAI221_X1 port map( B1 => n11734, B2 => n363, C1 => n10998, C2 => 
                           n374, A => n15634, ZN => n15633);
   U14179 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_31_23_port, B1 => 
                           n396, B2 => REGISTERS_35_23_port, C1 => n407, C2 => 
                           REGISTERS_39_23_port, ZN => n15634);
   U14180 : OAI221_X1 port map( B1 => n11574, B2 => n418, C1 => n11702, C2 => 
                           n429, A => n15635, ZN => n15632);
   U14181 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_26_23_port, B1 => 
                           n451, B2 => REGISTERS_30_23_port, C1 => n462, C2 => 
                           REGISTERS_34_23_port, ZN => n15635);
   U14182 : OAI221_X1 port map( B1 => n11414, B2 => n473, C1 => n11542, C2 => 
                           n484, A => n15636, ZN => n15631);
   U14183 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_21_23_port, B1 => 
                           n506, B2 => REGISTERS_25_23_port, C1 => n517, C2 => 
                           REGISTERS_29_23_port, ZN => n15636);
   U14184 : OAI221_X1 port map( B1 => n11254, B2 => n528, C1 => n11382, C2 => 
                           n539, A => n15637, ZN => n15630);
   U14185 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_24_23_port, B1 => 
                           n561, B2 => REGISTERS_22_23_port, C1 => n572, C2 => 
                           REGISTERS_20_23_port, ZN => n15637);
   U14186 : AOI22_X1 port map( A1 => n13880, A2 => n5104, B1 => n13881, B2 => 
                           n5105, ZN => n15598);
   U14187 : NOR4_X1 port map( A1 => n15640, A2 => n15641, A3 => n15642, A4 => 
                           n15643, ZN => n15639);
   U14188 : OAI221_X1 port map( B1 => n11062, B2 => n308, C1 => n10998, C2 => 
                           n319, A => n15644, ZN => n15643);
   U14189 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_14_23_port, B1 => 
                           n13808, B2 => REGISTERS_38_23_port, C1 => n13889, C2
                           => REGISTERS_39_23_port, ZN => n15644);
   U14190 : OAI221_X1 port map( B1 => n10902, B2 => n13810, C1 => n10838, C2 =>
                           n13890, A => n15645, ZN => n15642);
   U14191 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_23_port, B1 => 
                           n345, B2 => REGISTERS_9_23_port, C1 => n13812, C2 =>
                           REGISTERS_16_23_port, ZN => n15645);
   U14192 : OAI221_X1 port map( B1 => n10742, B2 => n303, C1 => n10678, C2 => 
                           n13893, A => n15646, ZN => n15641);
   U14193 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_23_port, B1 => 
                           n356, B2 => REGISTERS_4_23_port, C1 => n13818, C2 =>
                           REGISTERS_11_23_port, ZN => n15646);
   U14194 : OAI221_X1 port map( B1 => n11606, B2 => n304, C1 => n10550, C2 => 
                           n13896, A => n15647, ZN => n15640);
   U14195 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_23_port, B1 => 
                           n13826, B2 => REGISTERS_0_23_port, C1 => n13824, C2 
                           => REGISTERS_6_23_port, ZN => n15647);
   U14196 : NOR4_X1 port map( A1 => n15648, A2 => n15649, A3 => n15650, A4 => 
                           n15651, ZN => n15638);
   U14197 : OAI221_X1 port map( B1 => n11670, B2 => n363, C1 => n10934, C2 => 
                           n374, A => n15652, ZN => n15651);
   U14198 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_29_23_port, B1 => 
                           n396, B2 => REGISTERS_33_23_port, C1 => n407, C2 => 
                           REGISTERS_37_23_port, ZN => n15652);
   U14199 : OAI221_X1 port map( B1 => n11510, B2 => n418, C1 => n11638, C2 => 
                           n429, A => n15653, ZN => n15650);
   U14200 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_24_23_port, B1 => 
                           n451, B2 => REGISTERS_28_23_port, C1 => n462, C2 => 
                           REGISTERS_32_23_port, ZN => n15653);
   U14201 : OAI221_X1 port map( B1 => n11350, B2 => n473, C1 => n11478, C2 => 
                           n484, A => n15654, ZN => n15649);
   U14202 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_19_23_port, B1 => 
                           n506, B2 => REGISTERS_23_23_port, C1 => n517, C2 => 
                           REGISTERS_27_23_port, ZN => n15654);
   U14203 : OAI221_X1 port map( B1 => n11190, B2 => n528, C1 => n11318, C2 => 
                           n539, A => n15655, ZN => n15648);
   U14204 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_22_23_port, B1 => 
                           n561, B2 => REGISTERS_20_23_port, C1 => n572, C2 => 
                           REGISTERS_18_23_port, ZN => n15655);
   U14205 : NOR4_X1 port map( A1 => n15658, A2 => n15659, A3 => n15660, A4 => 
                           n15661, ZN => n15657);
   U14206 : OAI221_X1 port map( B1 => n11030, B2 => n308, C1 => n10966, C2 => 
                           n319, A => n15662, ZN => n15661);
   U14207 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_13_23_port, B1 => 
                           n13808, B2 => REGISTERS_37_23_port, C1 => n13889, C2
                           => REGISTERS_38_23_port, ZN => n15662);
   U14208 : OAI221_X1 port map( B1 => n10870, B2 => n13810, C1 => n10806, C2 =>
                           n13890, A => n15663, ZN => n15660);
   U14209 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_23_port, B1 => 
                           n345, B2 => REGISTERS_8_23_port, C1 => n13812, C2 =>
                           REGISTERS_15_23_port, ZN => n15663);
   U14210 : OAI221_X1 port map( B1 => n10710, B2 => n303, C1 => n10646, C2 => 
                           n13893, A => n15664, ZN => n15659);
   U14211 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_23_port, B1 => 
                           n356, B2 => REGISTERS_3_23_port, C1 => n13818, C2 =>
                           REGISTERS_10_23_port, ZN => n15664);
   U14212 : OAI221_X1 port map( B1 => n11574, B2 => n304, C1 => n10472, C2 => 
                           n13896, A => n15665, ZN => n15658);
   U14213 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_23_port, B1 => 
                           n13917, B2 => REGISTERS_39_23_port, C1 => n13824, C2
                           => REGISTERS_5_23_port, ZN => n15665);
   U14214 : NOR4_X1 port map( A1 => n15666, A2 => n15667, A3 => n15668, A4 => 
                           n15669, ZN => n15656);
   U14215 : OAI221_X1 port map( B1 => n11638, B2 => n363, C1 => n10902, C2 => 
                           n374, A => n15670, ZN => n15669);
   U14216 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_28_23_port, B1 => 
                           n396, B2 => REGISTERS_32_23_port, C1 => n407, C2 => 
                           REGISTERS_36_23_port, ZN => n15670);
   U14217 : OAI221_X1 port map( B1 => n11478, B2 => n418, C1 => n11606, C2 => 
                           n429, A => n15671, ZN => n15668);
   U14218 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_23_23_port, B1 => 
                           n451, B2 => REGISTERS_27_23_port, C1 => n462, C2 => 
                           REGISTERS_31_23_port, ZN => n15671);
   U14219 : OAI221_X1 port map( B1 => n11318, B2 => n473, C1 => n11446, C2 => 
                           n484, A => n15672, ZN => n15667);
   U14220 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_18_23_port, B1 => 
                           n506, B2 => REGISTERS_22_23_port, C1 => n517, C2 => 
                           REGISTERS_26_23_port, ZN => n15672);
   U14221 : OAI221_X1 port map( B1 => n11158, B2 => n528, C1 => n11286, C2 => 
                           n539, A => n15673, ZN => n15666);
   U14222 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_21_23_port, B1 => 
                           n561, B2 => REGISTERS_19_23_port, C1 => n572, C2 => 
                           REGISTERS_17_23_port, ZN => n15673);
   U14223 : NAND3_X1 port map( A1 => n15674, A2 => n15675, A3 => n15676, ZN => 
                           n11880);
   U14224 : AOI221_X1 port map( B1 => n13792, B2 => n5109, C1 => n13793, C2 => 
                           MEM_IN(24), A => n15677, ZN => n15676);
   U14225 : OAI22_X1 port map( A1 => n10469, A2 => n251, B1 => n5111, B2 => 
                           n121, ZN => n15677);
   U14226 : NOR2_X1 port map( A1 => n5704, A2 => n13796, ZN => n5702);
   U14227 : INV_X1 port map( A => MEM_IN(24), ZN => n5704);
   U14228 : AOI22_X1 port map( A1 => n197, A2 => n5112, B1 => n150, B2 => n5113
                           , ZN => n15675);
   U14229 : NOR4_X1 port map( A1 => n15680, A2 => n15681, A3 => n15682, A4 => 
                           n15683, ZN => n15679);
   U14230 : OAI221_X1 port map( B1 => n11093, B2 => n308, C1 => n11029, C2 => 
                           n319, A => n15684, ZN => n15683);
   U14231 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_15_24_port, B1 => 
                           n13807, B2 => REGISTERS_11_24_port, C1 => n13808, C2
                           => REGISTERS_39_24_port, ZN => n15684);
   U14232 : OAI221_X1 port map( B1 => n10805, B2 => n13809, C1 => n10933, C2 =>
                           n13810, A => n15685, ZN => n15682);
   U14233 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_24_port, B1 =>
                           n13813, B2 => REGISTERS_6_24_port, C1 => n349, C2 =>
                           REGISTERS_10_24_port, ZN => n15685);
   U14234 : OAI221_X1 port map( B1 => n10645, B2 => n13815, C1 => n10773, C2 =>
                           n303, A => n15686, ZN => n15681);
   U14235 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_24_port, B1 =>
                           n13819, B2 => REGISTERS_2_24_port, C1 => n360, C2 =>
                           REGISTERS_5_24_port, ZN => n15686);
   U14236 : OAI221_X1 port map( B1 => n10613, B2 => n13821, C1 => n11637, C2 =>
                           n304, A => n15687, ZN => n15680);
   U14237 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_24_port, B1 => 
                           n13825, B2 => REGISTERS_0_24_port, C1 => n13826, C2 
                           => REGISTERS_1_24_port, ZN => n15687);
   U14238 : NOR4_X1 port map( A1 => n15688, A2 => n15689, A3 => n15690, A4 => 
                           n15691, ZN => n15678);
   U14239 : OAI221_X1 port map( B1 => n11701, B2 => n363, C1 => n10965, C2 => 
                           n374, A => n15692, ZN => n15691);
   U14240 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_30_24_port, B1 => 
                           n396, B2 => REGISTERS_34_24_port, C1 => n407, C2 => 
                           REGISTERS_38_24_port, ZN => n15692);
   U14241 : OAI221_X1 port map( B1 => n11541, B2 => n418, C1 => n11669, C2 => 
                           n429, A => n15693, ZN => n15690);
   U14242 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_25_24_port, B1 => 
                           n451, B2 => REGISTERS_29_24_port, C1 => n462, C2 => 
                           REGISTERS_33_24_port, ZN => n15693);
   U14243 : OAI221_X1 port map( B1 => n11381, B2 => n473, C1 => n11509, C2 => 
                           n484, A => n15694, ZN => n15689);
   U14244 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_20_24_port, B1 => 
                           n506, B2 => REGISTERS_24_24_port, C1 => n517, C2 => 
                           REGISTERS_28_24_port, ZN => n15694);
   U14245 : OAI221_X1 port map( B1 => n11221, B2 => n528, C1 => n11349, C2 => 
                           n539, A => n15695, ZN => n15688);
   U14246 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_23_24_port, B1 => 
                           n561, B2 => REGISTERS_21_24_port, C1 => n572, C2 => 
                           REGISTERS_19_24_port, ZN => n15695);
   U14247 : NOR4_X1 port map( A1 => n15698, A2 => n15699, A3 => n15700, A4 => 
                           n15701, ZN => n15697);
   U14248 : OAI221_X1 port map( B1 => n11125, B2 => n308, C1 => n11061, C2 => 
                           n319, A => n15702, ZN => n15701);
   U14249 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_16_24_port, B1 => 
                           n119, B2 => REGISTERS_14_24_port, C1 => n13807, C2 
                           => REGISTERS_12_24_port, ZN => n15702);
   U14250 : OAI221_X1 port map( B1 => n11093, B2 => n13863, C1 => n10837, C2 =>
                           n13809, A => n15703, ZN => n15700);
   U14251 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_24_port, B1 => 
                           n13865, B2 => REGISTERS_9_24_port, C1 => n13813, C2 
                           => REGISTERS_7_24_port, ZN => n15703);
   U14252 : OAI221_X1 port map( B1 => n10933, B2 => n13866, C1 => n10677, C2 =>
                           n13815, A => n15704, ZN => n15699);
   U14253 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_24_port, B1 => 
                           n13868, B2 => REGISTERS_36_24_port, C1 => n13819, C2
                           => REGISTERS_3_24_port, ZN => n15704);
   U14254 : OAI221_X1 port map( B1 => n10773, B2 => n13869, C1 => n10645, C2 =>
                           n13821, A => n15705, ZN => n15698);
   U14255 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_24_port, B1 => 
                           n13871, B2 => REGISTERS_0_24_port, C1 => n13825, C2 
                           => REGISTERS_1_24_port, ZN => n15705);
   U14256 : NOR4_X1 port map( A1 => n15706, A2 => n15707, A3 => n15708, A4 => 
                           n15709, ZN => n15696);
   U14257 : OAI221_X1 port map( B1 => n11733, B2 => n363, C1 => n10997, C2 => 
                           n374, A => n15710, ZN => n15709);
   U14258 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_31_24_port, B1 => 
                           n396, B2 => REGISTERS_35_24_port, C1 => n407, C2 => 
                           REGISTERS_39_24_port, ZN => n15710);
   U14259 : OAI221_X1 port map( B1 => n11573, B2 => n418, C1 => n11701, C2 => 
                           n429, A => n15711, ZN => n15708);
   U14260 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_26_24_port, B1 => 
                           n451, B2 => REGISTERS_30_24_port, C1 => n462, C2 => 
                           REGISTERS_34_24_port, ZN => n15711);
   U14261 : OAI221_X1 port map( B1 => n11413, B2 => n473, C1 => n11541, C2 => 
                           n484, A => n15712, ZN => n15707);
   U14262 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_21_24_port, B1 => 
                           n506, B2 => REGISTERS_25_24_port, C1 => n517, C2 => 
                           REGISTERS_29_24_port, ZN => n15712);
   U14263 : OAI221_X1 port map( B1 => n11253, B2 => n528, C1 => n11381, C2 => 
                           n539, A => n15713, ZN => n15706);
   U14264 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_24_24_port, B1 => 
                           n561, B2 => REGISTERS_22_24_port, C1 => n572, C2 => 
                           REGISTERS_20_24_port, ZN => n15713);
   U14265 : AOI22_X1 port map( A1 => n13880, A2 => n5114, B1 => n13881, B2 => 
                           n5115, ZN => n15674);
   U14266 : NOR4_X1 port map( A1 => n15716, A2 => n15717, A3 => n15718, A4 => 
                           n15719, ZN => n15715);
   U14267 : OAI221_X1 port map( B1 => n11061, B2 => n308, C1 => n10997, C2 => 
                           n319, A => n15720, ZN => n15719);
   U14268 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_14_24_port, B1 => 
                           n13808, B2 => REGISTERS_38_24_port, C1 => n13889, C2
                           => REGISTERS_39_24_port, ZN => n15720);
   U14269 : OAI221_X1 port map( B1 => n10901, B2 => n13810, C1 => n10837, C2 =>
                           n13890, A => n15721, ZN => n15718);
   U14270 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_24_port, B1 => 
                           n345, B2 => REGISTERS_9_24_port, C1 => n13812, C2 =>
                           REGISTERS_16_24_port, ZN => n15721);
   U14271 : OAI221_X1 port map( B1 => n10741, B2 => n303, C1 => n10677, C2 => 
                           n13893, A => n15722, ZN => n15717);
   U14272 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_24_port, B1 => 
                           n356, B2 => REGISTERS_4_24_port, C1 => n13818, C2 =>
                           REGISTERS_11_24_port, ZN => n15722);
   U14273 : OAI221_X1 port map( B1 => n11605, B2 => n304, C1 => n10549, C2 => 
                           n13896, A => n15723, ZN => n15716);
   U14274 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_24_port, B1 => 
                           n13826, B2 => REGISTERS_0_24_port, C1 => n13824, C2 
                           => REGISTERS_6_24_port, ZN => n15723);
   U14275 : NOR4_X1 port map( A1 => n15724, A2 => n15725, A3 => n15726, A4 => 
                           n15727, ZN => n15714);
   U14276 : OAI221_X1 port map( B1 => n11669, B2 => n363, C1 => n10933, C2 => 
                           n374, A => n15728, ZN => n15727);
   U14277 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_29_24_port, B1 => 
                           n396, B2 => REGISTERS_33_24_port, C1 => n407, C2 => 
                           REGISTERS_37_24_port, ZN => n15728);
   U14278 : OAI221_X1 port map( B1 => n11509, B2 => n418, C1 => n11637, C2 => 
                           n429, A => n15729, ZN => n15726);
   U14279 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_24_24_port, B1 => 
                           n451, B2 => REGISTERS_28_24_port, C1 => n462, C2 => 
                           REGISTERS_32_24_port, ZN => n15729);
   U14280 : OAI221_X1 port map( B1 => n11349, B2 => n473, C1 => n11477, C2 => 
                           n484, A => n15730, ZN => n15725);
   U14281 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_19_24_port, B1 => 
                           n506, B2 => REGISTERS_23_24_port, C1 => n517, C2 => 
                           REGISTERS_27_24_port, ZN => n15730);
   U14282 : OAI221_X1 port map( B1 => n11189, B2 => n528, C1 => n11317, C2 => 
                           n539, A => n15731, ZN => n15724);
   U14283 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_22_24_port, B1 => 
                           n561, B2 => REGISTERS_20_24_port, C1 => n572, C2 => 
                           REGISTERS_18_24_port, ZN => n15731);
   U14284 : NOR4_X1 port map( A1 => n15734, A2 => n15735, A3 => n15736, A4 => 
                           n15737, ZN => n15733);
   U14285 : OAI221_X1 port map( B1 => n11029, B2 => n308, C1 => n10965, C2 => 
                           n319, A => n15738, ZN => n15737);
   U14286 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_13_24_port, B1 => 
                           n13808, B2 => REGISTERS_37_24_port, C1 => n13889, C2
                           => REGISTERS_38_24_port, ZN => n15738);
   U14287 : OAI221_X1 port map( B1 => n10869, B2 => n13810, C1 => n10805, C2 =>
                           n13890, A => n15739, ZN => n15736);
   U14288 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_24_port, B1 => 
                           n345, B2 => REGISTERS_8_24_port, C1 => n13812, C2 =>
                           REGISTERS_15_24_port, ZN => n15739);
   U14289 : OAI221_X1 port map( B1 => n10709, B2 => n303, C1 => n10645, C2 => 
                           n13893, A => n15740, ZN => n15735);
   U14290 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_24_port, B1 => 
                           n356, B2 => REGISTERS_3_24_port, C1 => n13818, C2 =>
                           REGISTERS_10_24_port, ZN => n15740);
   U14291 : OAI221_X1 port map( B1 => n11573, B2 => n304, C1 => n10469, C2 => 
                           n13896, A => n15741, ZN => n15734);
   U14292 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_24_port, B1 => 
                           n13917, B2 => REGISTERS_39_24_port, C1 => n13824, C2
                           => REGISTERS_5_24_port, ZN => n15741);
   U14293 : NOR4_X1 port map( A1 => n15742, A2 => n15743, A3 => n15744, A4 => 
                           n15745, ZN => n15732);
   U14294 : OAI221_X1 port map( B1 => n11637, B2 => n363, C1 => n10901, C2 => 
                           n374, A => n15746, ZN => n15745);
   U14295 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_28_24_port, B1 => 
                           n396, B2 => REGISTERS_32_24_port, C1 => n407, C2 => 
                           REGISTERS_36_24_port, ZN => n15746);
   U14296 : OAI221_X1 port map( B1 => n11477, B2 => n418, C1 => n11605, C2 => 
                           n429, A => n15747, ZN => n15744);
   U14297 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_23_24_port, B1 => 
                           n451, B2 => REGISTERS_27_24_port, C1 => n462, C2 => 
                           REGISTERS_31_24_port, ZN => n15747);
   U14298 : OAI221_X1 port map( B1 => n11317, B2 => n473, C1 => n11445, C2 => 
                           n484, A => n15748, ZN => n15743);
   U14299 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_18_24_port, B1 => 
                           n506, B2 => REGISTERS_22_24_port, C1 => n517, C2 => 
                           REGISTERS_26_24_port, ZN => n15748);
   U14300 : OAI221_X1 port map( B1 => n11157, B2 => n528, C1 => n11285, C2 => 
                           n539, A => n15749, ZN => n15742);
   U14301 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_21_24_port, B1 => 
                           n561, B2 => REGISTERS_19_24_port, C1 => n572, C2 => 
                           REGISTERS_17_24_port, ZN => n15749);
   U14302 : NAND3_X1 port map( A1 => n15750, A2 => n15751, A3 => n15752, ZN => 
                           n11879);
   U14303 : AOI221_X1 port map( B1 => n13792, B2 => n5119, C1 => n13793, C2 => 
                           MEM_IN(25), A => n15753, ZN => n15752);
   U14304 : OAI22_X1 port map( A1 => n10466, A2 => n251, B1 => n5121, B2 => 
                           n121, ZN => n15753);
   U14305 : NOR2_X1 port map( A1 => n5711, A2 => n13796, ZN => n5709);
   U14306 : INV_X1 port map( A => MEM_IN(25), ZN => n5711);
   U14307 : AOI22_X1 port map( A1 => n197, A2 => n5122, B1 => n150, B2 => n5123
                           , ZN => n15751);
   U14308 : NOR4_X1 port map( A1 => n15756, A2 => n15757, A3 => n15758, A4 => 
                           n15759, ZN => n15755);
   U14309 : OAI221_X1 port map( B1 => n11092, B2 => n308, C1 => n11028, C2 => 
                           n319, A => n15760, ZN => n15759);
   U14310 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_15_25_port, B1 => 
                           n13807, B2 => REGISTERS_11_25_port, C1 => n13808, C2
                           => REGISTERS_39_25_port, ZN => n15760);
   U14311 : OAI221_X1 port map( B1 => n10804, B2 => n13809, C1 => n10932, C2 =>
                           n13810, A => n15761, ZN => n15758);
   U14312 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_25_port, B1 =>
                           n13813, B2 => REGISTERS_6_25_port, C1 => n349, C2 =>
                           REGISTERS_10_25_port, ZN => n15761);
   U14313 : OAI221_X1 port map( B1 => n10644, B2 => n13815, C1 => n10772, C2 =>
                           n303, A => n15762, ZN => n15757);
   U14314 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_25_port, B1 =>
                           n13819, B2 => REGISTERS_2_25_port, C1 => n360, C2 =>
                           REGISTERS_5_25_port, ZN => n15762);
   U14315 : OAI221_X1 port map( B1 => n10612, B2 => n13821, C1 => n11636, C2 =>
                           n304, A => n15763, ZN => n15756);
   U14316 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_25_port, B1 => 
                           n13825, B2 => REGISTERS_0_25_port, C1 => n13826, C2 
                           => REGISTERS_1_25_port, ZN => n15763);
   U14317 : NOR4_X1 port map( A1 => n15764, A2 => n15765, A3 => n15766, A4 => 
                           n15767, ZN => n15754);
   U14318 : OAI221_X1 port map( B1 => n11700, B2 => n363, C1 => n10964, C2 => 
                           n374, A => n15768, ZN => n15767);
   U14319 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_30_25_port, B1 => 
                           n396, B2 => REGISTERS_34_25_port, C1 => n407, C2 => 
                           REGISTERS_38_25_port, ZN => n15768);
   U14320 : OAI221_X1 port map( B1 => n11540, B2 => n418, C1 => n11668, C2 => 
                           n429, A => n15769, ZN => n15766);
   U14321 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_25_25_port, B1 => 
                           n451, B2 => REGISTERS_29_25_port, C1 => n462, C2 => 
                           REGISTERS_33_25_port, ZN => n15769);
   U14322 : OAI221_X1 port map( B1 => n11380, B2 => n473, C1 => n11508, C2 => 
                           n484, A => n15770, ZN => n15765);
   U14323 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_20_25_port, B1 => 
                           n506, B2 => REGISTERS_24_25_port, C1 => n517, C2 => 
                           REGISTERS_28_25_port, ZN => n15770);
   U14324 : OAI221_X1 port map( B1 => n11220, B2 => n528, C1 => n11348, C2 => 
                           n539, A => n15771, ZN => n15764);
   U14325 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_23_25_port, B1 => 
                           n561, B2 => REGISTERS_21_25_port, C1 => n572, C2 => 
                           REGISTERS_19_25_port, ZN => n15771);
   U14326 : NOR4_X1 port map( A1 => n15774, A2 => n15775, A3 => n15776, A4 => 
                           n15777, ZN => n15773);
   U14327 : OAI221_X1 port map( B1 => n11124, B2 => n308, C1 => n11060, C2 => 
                           n319, A => n15778, ZN => n15777);
   U14328 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_16_25_port, B1 => 
                           n119, B2 => REGISTERS_14_25_port, C1 => n13807, C2 
                           => REGISTERS_12_25_port, ZN => n15778);
   U14329 : OAI221_X1 port map( B1 => n11092, B2 => n13863, C1 => n10836, C2 =>
                           n13809, A => n15779, ZN => n15776);
   U14330 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_25_port, B1 => 
                           n13865, B2 => REGISTERS_9_25_port, C1 => n13813, C2 
                           => REGISTERS_7_25_port, ZN => n15779);
   U14331 : OAI221_X1 port map( B1 => n10932, B2 => n13866, C1 => n10676, C2 =>
                           n13815, A => n15780, ZN => n15775);
   U14332 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_25_port, B1 => 
                           n13868, B2 => REGISTERS_36_25_port, C1 => n13819, C2
                           => REGISTERS_3_25_port, ZN => n15780);
   U14333 : OAI221_X1 port map( B1 => n10772, B2 => n13869, C1 => n10644, C2 =>
                           n13821, A => n15781, ZN => n15774);
   U14334 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_25_port, B1 => 
                           n13871, B2 => REGISTERS_0_25_port, C1 => n13825, C2 
                           => REGISTERS_1_25_port, ZN => n15781);
   U14335 : NOR4_X1 port map( A1 => n15782, A2 => n15783, A3 => n15784, A4 => 
                           n15785, ZN => n15772);
   U14336 : OAI221_X1 port map( B1 => n11732, B2 => n363, C1 => n10996, C2 => 
                           n374, A => n15786, ZN => n15785);
   U14337 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_31_25_port, B1 => 
                           n396, B2 => REGISTERS_35_25_port, C1 => n407, C2 => 
                           REGISTERS_39_25_port, ZN => n15786);
   U14338 : OAI221_X1 port map( B1 => n11572, B2 => n418, C1 => n11700, C2 => 
                           n429, A => n15787, ZN => n15784);
   U14339 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_26_25_port, B1 => 
                           n451, B2 => REGISTERS_30_25_port, C1 => n462, C2 => 
                           REGISTERS_34_25_port, ZN => n15787);
   U14340 : OAI221_X1 port map( B1 => n11412, B2 => n473, C1 => n11540, C2 => 
                           n484, A => n15788, ZN => n15783);
   U14341 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_21_25_port, B1 => 
                           n506, B2 => REGISTERS_25_25_port, C1 => n517, C2 => 
                           REGISTERS_29_25_port, ZN => n15788);
   U14342 : OAI221_X1 port map( B1 => n11252, B2 => n528, C1 => n11380, C2 => 
                           n539, A => n15789, ZN => n15782);
   U14343 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_24_25_port, B1 => 
                           n561, B2 => REGISTERS_22_25_port, C1 => n572, C2 => 
                           REGISTERS_20_25_port, ZN => n15789);
   U14344 : AOI22_X1 port map( A1 => n13880, A2 => n5124, B1 => n13881, B2 => 
                           n5125, ZN => n15750);
   U14345 : NOR4_X1 port map( A1 => n15792, A2 => n15793, A3 => n15794, A4 => 
                           n15795, ZN => n15791);
   U14346 : OAI221_X1 port map( B1 => n11060, B2 => n308, C1 => n10996, C2 => 
                           n319, A => n15796, ZN => n15795);
   U14347 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_14_25_port, B1 => 
                           n13808, B2 => REGISTERS_38_25_port, C1 => n13889, C2
                           => REGISTERS_39_25_port, ZN => n15796);
   U14348 : OAI221_X1 port map( B1 => n10900, B2 => n13810, C1 => n10836, C2 =>
                           n13890, A => n15797, ZN => n15794);
   U14349 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_25_port, B1 => 
                           n345, B2 => REGISTERS_9_25_port, C1 => n13812, C2 =>
                           REGISTERS_16_25_port, ZN => n15797);
   U14350 : OAI221_X1 port map( B1 => n10740, B2 => n303, C1 => n10676, C2 => 
                           n13893, A => n15798, ZN => n15793);
   U14351 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_25_port, B1 => 
                           n356, B2 => REGISTERS_4_25_port, C1 => n13818, C2 =>
                           REGISTERS_11_25_port, ZN => n15798);
   U14352 : OAI221_X1 port map( B1 => n11604, B2 => n304, C1 => n10548, C2 => 
                           n13896, A => n15799, ZN => n15792);
   U14353 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_25_port, B1 => 
                           n13826, B2 => REGISTERS_0_25_port, C1 => n13824, C2 
                           => REGISTERS_6_25_port, ZN => n15799);
   U14354 : NOR4_X1 port map( A1 => n15800, A2 => n15801, A3 => n15802, A4 => 
                           n15803, ZN => n15790);
   U14355 : OAI221_X1 port map( B1 => n11668, B2 => n363, C1 => n10932, C2 => 
                           n374, A => n15804, ZN => n15803);
   U14356 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_29_25_port, B1 => 
                           n396, B2 => REGISTERS_33_25_port, C1 => n407, C2 => 
                           REGISTERS_37_25_port, ZN => n15804);
   U14357 : OAI221_X1 port map( B1 => n11508, B2 => n418, C1 => n11636, C2 => 
                           n429, A => n15805, ZN => n15802);
   U14358 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_24_25_port, B1 => 
                           n451, B2 => REGISTERS_28_25_port, C1 => n462, C2 => 
                           REGISTERS_32_25_port, ZN => n15805);
   U14359 : OAI221_X1 port map( B1 => n11348, B2 => n473, C1 => n11476, C2 => 
                           n484, A => n15806, ZN => n15801);
   U14360 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_19_25_port, B1 => 
                           n506, B2 => REGISTERS_23_25_port, C1 => n517, C2 => 
                           REGISTERS_27_25_port, ZN => n15806);
   U14361 : OAI221_X1 port map( B1 => n11188, B2 => n528, C1 => n11316, C2 => 
                           n539, A => n15807, ZN => n15800);
   U14362 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_22_25_port, B1 => 
                           n561, B2 => REGISTERS_20_25_port, C1 => n572, C2 => 
                           REGISTERS_18_25_port, ZN => n15807);
   U14363 : NOR4_X1 port map( A1 => n15810, A2 => n15811, A3 => n15812, A4 => 
                           n15813, ZN => n15809);
   U14364 : OAI221_X1 port map( B1 => n11028, B2 => n308, C1 => n10964, C2 => 
                           n319, A => n15814, ZN => n15813);
   U14365 : AOI222_X1 port map( A1 => n330, A2 => REGISTERS_13_25_port, B1 => 
                           n13808, B2 => REGISTERS_37_25_port, C1 => n13889, C2
                           => REGISTERS_38_25_port, ZN => n15814);
   U14366 : OAI221_X1 port map( B1 => n10868, B2 => n13810, C1 => n10804, C2 =>
                           n13890, A => n15815, ZN => n15812);
   U14367 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_25_port, B1 => 
                           n345, B2 => REGISTERS_8_25_port, C1 => n13812, C2 =>
                           REGISTERS_15_25_port, ZN => n15815);
   U14368 : OAI221_X1 port map( B1 => n10708, B2 => n303, C1 => n10644, C2 => 
                           n13893, A => n15816, ZN => n15811);
   U14369 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_25_port, B1 => 
                           n356, B2 => REGISTERS_3_25_port, C1 => n13818, C2 =>
                           REGISTERS_10_25_port, ZN => n15816);
   U14370 : OAI221_X1 port map( B1 => n11572, B2 => n304, C1 => n10466, C2 => 
                           n13896, A => n15817, ZN => n15810);
   U14371 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_25_port, B1 => 
                           n13917, B2 => REGISTERS_39_25_port, C1 => n13824, C2
                           => REGISTERS_5_25_port, ZN => n15817);
   U14372 : NOR4_X1 port map( A1 => n15818, A2 => n15819, A3 => n15820, A4 => 
                           n15821, ZN => n15808);
   U14373 : OAI221_X1 port map( B1 => n11636, B2 => n363, C1 => n10900, C2 => 
                           n374, A => n15822, ZN => n15821);
   U14374 : AOI222_X1 port map( A1 => n385, A2 => REGISTERS_28_25_port, B1 => 
                           n396, B2 => REGISTERS_32_25_port, C1 => n407, C2 => 
                           REGISTERS_36_25_port, ZN => n15822);
   U14375 : OAI221_X1 port map( B1 => n11476, B2 => n418, C1 => n11604, C2 => 
                           n429, A => n15823, ZN => n15820);
   U14376 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_23_25_port, B1 => 
                           n451, B2 => REGISTERS_27_25_port, C1 => n462, C2 => 
                           REGISTERS_31_25_port, ZN => n15823);
   U14377 : OAI221_X1 port map( B1 => n11316, B2 => n473, C1 => n11444, C2 => 
                           n484, A => n15824, ZN => n15819);
   U14378 : AOI222_X1 port map( A1 => n495, A2 => REGISTERS_18_25_port, B1 => 
                           n506, B2 => REGISTERS_22_25_port, C1 => n517, C2 => 
                           REGISTERS_26_25_port, ZN => n15824);
   U14379 : OAI221_X1 port map( B1 => n11156, B2 => n528, C1 => n11284, C2 => 
                           n539, A => n15825, ZN => n15818);
   U14380 : AOI222_X1 port map( A1 => n550, A2 => REGISTERS_21_25_port, B1 => 
                           n561, B2 => REGISTERS_19_25_port, C1 => n572, C2 => 
                           REGISTERS_17_25_port, ZN => n15825);
   U14381 : NAND3_X1 port map( A1 => n15826, A2 => n15827, A3 => n15828, ZN => 
                           n11878);
   U14382 : AOI221_X1 port map( B1 => n13792, B2 => n5129, C1 => n13793, C2 => 
                           MEM_IN(26), A => n15829, ZN => n15828);
   U14383 : OAI22_X1 port map( A1 => n10463, A2 => n251, B1 => n5131, B2 => 
                           n121, ZN => n15829);
   U14384 : NOR2_X1 port map( A1 => n5718, A2 => n13796, ZN => n5716);
   U14385 : INV_X1 port map( A => MEM_IN(26), ZN => n5718);
   U14386 : AOI22_X1 port map( A1 => n197, A2 => n5132, B1 => n150, B2 => n5133
                           , ZN => n15827);
   U14387 : NOR4_X1 port map( A1 => n15832, A2 => n15833, A3 => n15834, A4 => 
                           n15835, ZN => n15831);
   U14388 : OAI221_X1 port map( B1 => n11091, B2 => n307, C1 => n11027, C2 => 
                           n318, A => n15836, ZN => n15835);
   U14389 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_15_26_port, B1 => 
                           n13807, B2 => REGISTERS_11_26_port, C1 => n13808, C2
                           => REGISTERS_39_26_port, ZN => n15836);
   U14390 : OAI221_X1 port map( B1 => n10803, B2 => n13809, C1 => n10931, C2 =>
                           n13810, A => n15837, ZN => n15834);
   U14391 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_26_port, B1 =>
                           n13813, B2 => REGISTERS_6_26_port, C1 => n349, C2 =>
                           REGISTERS_10_26_port, ZN => n15837);
   U14392 : OAI221_X1 port map( B1 => n10643, B2 => n13815, C1 => n10771, C2 =>
                           n303, A => n15838, ZN => n15833);
   U14393 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_26_port, B1 =>
                           n13819, B2 => REGISTERS_2_26_port, C1 => n360, C2 =>
                           REGISTERS_5_26_port, ZN => n15838);
   U14394 : OAI221_X1 port map( B1 => n10611, B2 => n13821, C1 => n11635, C2 =>
                           n304, A => n15839, ZN => n15832);
   U14395 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_26_port, B1 => 
                           n13825, B2 => REGISTERS_0_26_port, C1 => n13826, C2 
                           => REGISTERS_1_26_port, ZN => n15839);
   U14396 : NOR4_X1 port map( A1 => n15840, A2 => n15841, A3 => n15842, A4 => 
                           n15843, ZN => n15830);
   U14397 : OAI221_X1 port map( B1 => n11699, B2 => n362, C1 => n10963, C2 => 
                           n374, A => n15844, ZN => n15843);
   U14398 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_30_26_port, B1 => 
                           n395, B2 => REGISTERS_34_26_port, C1 => n406, C2 => 
                           REGISTERS_38_26_port, ZN => n15844);
   U14399 : OAI221_X1 port map( B1 => n11539, B2 => n417, C1 => n11667, C2 => 
                           n428, A => n15845, ZN => n15842);
   U14400 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_25_26_port, B1 => 
                           n450, B2 => REGISTERS_29_26_port, C1 => n461, C2 => 
                           REGISTERS_33_26_port, ZN => n15845);
   U14401 : OAI221_X1 port map( B1 => n11379, B2 => n472, C1 => n11507, C2 => 
                           n483, A => n15846, ZN => n15841);
   U14402 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_20_26_port, B1 => 
                           n505, B2 => REGISTERS_24_26_port, C1 => n516, C2 => 
                           REGISTERS_28_26_port, ZN => n15846);
   U14403 : OAI221_X1 port map( B1 => n11219, B2 => n527, C1 => n11347, C2 => 
                           n538, A => n15847, ZN => n15840);
   U14404 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_23_26_port, B1 => 
                           n560, B2 => REGISTERS_21_26_port, C1 => n571, C2 => 
                           REGISTERS_19_26_port, ZN => n15847);
   U14405 : NOR4_X1 port map( A1 => n15850, A2 => n15851, A3 => n15852, A4 => 
                           n15853, ZN => n15849);
   U14406 : OAI221_X1 port map( B1 => n11123, B2 => n307, C1 => n11059, C2 => 
                           n318, A => n15854, ZN => n15853);
   U14407 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_16_26_port, B1 => 
                           n119, B2 => REGISTERS_14_26_port, C1 => n13807, C2 
                           => REGISTERS_12_26_port, ZN => n15854);
   U14408 : OAI221_X1 port map( B1 => n11091, B2 => n13863, C1 => n10835, C2 =>
                           n13809, A => n15855, ZN => n15852);
   U14409 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_26_port, B1 => 
                           n13865, B2 => REGISTERS_9_26_port, C1 => n13813, C2 
                           => REGISTERS_7_26_port, ZN => n15855);
   U14410 : OAI221_X1 port map( B1 => n10931, B2 => n13866, C1 => n10675, C2 =>
                           n13815, A => n15856, ZN => n15851);
   U14411 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_26_port, B1 => 
                           n13868, B2 => REGISTERS_36_26_port, C1 => n13819, C2
                           => REGISTERS_3_26_port, ZN => n15856);
   U14412 : OAI221_X1 port map( B1 => n10771, B2 => n13869, C1 => n10643, C2 =>
                           n13821, A => n15857, ZN => n15850);
   U14413 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_26_port, B1 => 
                           n13871, B2 => REGISTERS_0_26_port, C1 => n13825, C2 
                           => REGISTERS_1_26_port, ZN => n15857);
   U14414 : NOR4_X1 port map( A1 => n15858, A2 => n15859, A3 => n15860, A4 => 
                           n15861, ZN => n15848);
   U14415 : OAI221_X1 port map( B1 => n11731, B2 => n362, C1 => n10995, C2 => 
                           n373, A => n15862, ZN => n15861);
   U14416 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_31_26_port, B1 => 
                           n395, B2 => REGISTERS_35_26_port, C1 => n406, C2 => 
                           REGISTERS_39_26_port, ZN => n15862);
   U14417 : OAI221_X1 port map( B1 => n11571, B2 => n417, C1 => n11699, C2 => 
                           n428, A => n15863, ZN => n15860);
   U14418 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_26_26_port, B1 => 
                           n450, B2 => REGISTERS_30_26_port, C1 => n461, C2 => 
                           REGISTERS_34_26_port, ZN => n15863);
   U14419 : OAI221_X1 port map( B1 => n11411, B2 => n472, C1 => n11539, C2 => 
                           n483, A => n15864, ZN => n15859);
   U14420 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_21_26_port, B1 => 
                           n505, B2 => REGISTERS_25_26_port, C1 => n516, C2 => 
                           REGISTERS_29_26_port, ZN => n15864);
   U14421 : OAI221_X1 port map( B1 => n11251, B2 => n527, C1 => n11379, C2 => 
                           n538, A => n15865, ZN => n15858);
   U14422 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_24_26_port, B1 => 
                           n560, B2 => REGISTERS_22_26_port, C1 => n571, C2 => 
                           REGISTERS_20_26_port, ZN => n15865);
   U14423 : AOI22_X1 port map( A1 => n13880, A2 => n5134, B1 => n13881, B2 => 
                           n5135, ZN => n15826);
   U14424 : NOR4_X1 port map( A1 => n15868, A2 => n15869, A3 => n15870, A4 => 
                           n15871, ZN => n15867);
   U14425 : OAI221_X1 port map( B1 => n11059, B2 => n307, C1 => n10995, C2 => 
                           n318, A => n15872, ZN => n15871);
   U14426 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_14_26_port, B1 => 
                           n13808, B2 => REGISTERS_38_26_port, C1 => n13889, C2
                           => REGISTERS_39_26_port, ZN => n15872);
   U14427 : OAI221_X1 port map( B1 => n10899, B2 => n13810, C1 => n10835, C2 =>
                           n13890, A => n15873, ZN => n15870);
   U14428 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_26_port, B1 => 
                           n346, B2 => REGISTERS_9_26_port, C1 => n13812, C2 =>
                           REGISTERS_16_26_port, ZN => n15873);
   U14429 : OAI221_X1 port map( B1 => n10739, B2 => n303, C1 => n10675, C2 => 
                           n13893, A => n15874, ZN => n15869);
   U14430 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_26_port, B1 => 
                           n357, B2 => REGISTERS_4_26_port, C1 => n13818, C2 =>
                           REGISTERS_11_26_port, ZN => n15874);
   U14431 : OAI221_X1 port map( B1 => n11603, B2 => n304, C1 => n10547, C2 => 
                           n13896, A => n15875, ZN => n15868);
   U14432 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_26_port, B1 => 
                           n13826, B2 => REGISTERS_0_26_port, C1 => n13824, C2 
                           => REGISTERS_6_26_port, ZN => n15875);
   U14433 : NOR4_X1 port map( A1 => n15876, A2 => n15877, A3 => n15878, A4 => 
                           n15879, ZN => n15866);
   U14434 : OAI221_X1 port map( B1 => n11667, B2 => n362, C1 => n10931, C2 => 
                           n373, A => n15880, ZN => n15879);
   U14435 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_29_26_port, B1 => 
                           n395, B2 => REGISTERS_33_26_port, C1 => n406, C2 => 
                           REGISTERS_37_26_port, ZN => n15880);
   U14436 : OAI221_X1 port map( B1 => n11507, B2 => n417, C1 => n11635, C2 => 
                           n428, A => n15881, ZN => n15878);
   U14437 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_24_26_port, B1 => 
                           n450, B2 => REGISTERS_28_26_port, C1 => n461, C2 => 
                           REGISTERS_32_26_port, ZN => n15881);
   U14438 : OAI221_X1 port map( B1 => n11347, B2 => n472, C1 => n11475, C2 => 
                           n483, A => n15882, ZN => n15877);
   U14439 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_19_26_port, B1 => 
                           n505, B2 => REGISTERS_23_26_port, C1 => n516, C2 => 
                           REGISTERS_27_26_port, ZN => n15882);
   U14440 : OAI221_X1 port map( B1 => n11187, B2 => n527, C1 => n11315, C2 => 
                           n538, A => n15883, ZN => n15876);
   U14441 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_22_26_port, B1 => 
                           n560, B2 => REGISTERS_20_26_port, C1 => n571, C2 => 
                           REGISTERS_18_26_port, ZN => n15883);
   U14442 : NOR4_X1 port map( A1 => n15886, A2 => n15887, A3 => n15888, A4 => 
                           n15889, ZN => n15885);
   U14443 : OAI221_X1 port map( B1 => n11027, B2 => n307, C1 => n10963, C2 => 
                           n318, A => n15890, ZN => n15889);
   U14444 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_13_26_port, B1 => 
                           n13808, B2 => REGISTERS_37_26_port, C1 => n13889, C2
                           => REGISTERS_38_26_port, ZN => n15890);
   U14445 : OAI221_X1 port map( B1 => n10867, B2 => n13810, C1 => n10803, C2 =>
                           n13890, A => n15891, ZN => n15888);
   U14446 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_26_port, B1 => 
                           n346, B2 => REGISTERS_8_26_port, C1 => n13812, C2 =>
                           REGISTERS_15_26_port, ZN => n15891);
   U14447 : OAI221_X1 port map( B1 => n10707, B2 => n303, C1 => n10643, C2 => 
                           n13893, A => n15892, ZN => n15887);
   U14448 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_26_port, B1 => 
                           n357, B2 => REGISTERS_3_26_port, C1 => n13818, C2 =>
                           REGISTERS_10_26_port, ZN => n15892);
   U14449 : OAI221_X1 port map( B1 => n11571, B2 => n304, C1 => n10463, C2 => 
                           n13896, A => n15893, ZN => n15886);
   U14450 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_26_port, B1 => 
                           n13917, B2 => REGISTERS_39_26_port, C1 => n13824, C2
                           => REGISTERS_5_26_port, ZN => n15893);
   U14451 : NOR4_X1 port map( A1 => n15894, A2 => n15895, A3 => n15896, A4 => 
                           n15897, ZN => n15884);
   U14452 : OAI221_X1 port map( B1 => n11635, B2 => n362, C1 => n10899, C2 => 
                           n373, A => n15898, ZN => n15897);
   U14453 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_28_26_port, B1 => 
                           n395, B2 => REGISTERS_32_26_port, C1 => n406, C2 => 
                           REGISTERS_36_26_port, ZN => n15898);
   U14454 : OAI221_X1 port map( B1 => n11475, B2 => n417, C1 => n11603, C2 => 
                           n428, A => n15899, ZN => n15896);
   U14455 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_23_26_port, B1 => 
                           n450, B2 => REGISTERS_27_26_port, C1 => n461, C2 => 
                           REGISTERS_31_26_port, ZN => n15899);
   U14456 : OAI221_X1 port map( B1 => n11315, B2 => n472, C1 => n11443, C2 => 
                           n483, A => n15900, ZN => n15895);
   U14457 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_18_26_port, B1 => 
                           n505, B2 => REGISTERS_22_26_port, C1 => n516, C2 => 
                           REGISTERS_26_26_port, ZN => n15900);
   U14458 : OAI221_X1 port map( B1 => n11155, B2 => n527, C1 => n11283, C2 => 
                           n538, A => n15901, ZN => n15894);
   U14459 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_21_26_port, B1 => 
                           n560, B2 => REGISTERS_19_26_port, C1 => n571, C2 => 
                           REGISTERS_17_26_port, ZN => n15901);
   U14460 : NAND3_X1 port map( A1 => n15902, A2 => n15903, A3 => n15904, ZN => 
                           n11877);
   U14461 : AOI221_X1 port map( B1 => n13792, B2 => n5139, C1 => n13793, C2 => 
                           MEM_IN(27), A => n15905, ZN => n15904);
   U14462 : OAI22_X1 port map( A1 => n10460, A2 => n251, B1 => n5141, B2 => 
                           n121, ZN => n15905);
   U14463 : NOR2_X1 port map( A1 => n5725, A2 => n13796, ZN => n5723);
   U14464 : INV_X1 port map( A => MEM_IN(27), ZN => n5725);
   U14465 : AOI22_X1 port map( A1 => n197, A2 => n5142, B1 => n150, B2 => n5143
                           , ZN => n15903);
   U14466 : NOR4_X1 port map( A1 => n15908, A2 => n15909, A3 => n15910, A4 => 
                           n15911, ZN => n15907);
   U14467 : OAI221_X1 port map( B1 => n11090, B2 => n307, C1 => n11026, C2 => 
                           n318, A => n15912, ZN => n15911);
   U14468 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_15_27_port, B1 => 
                           n13807, B2 => REGISTERS_11_27_port, C1 => n13808, C2
                           => REGISTERS_39_27_port, ZN => n15912);
   U14469 : OAI221_X1 port map( B1 => n10802, B2 => n13809, C1 => n10930, C2 =>
                           n13810, A => n15913, ZN => n15910);
   U14470 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_27_port, B1 =>
                           n13813, B2 => REGISTERS_6_27_port, C1 => n349, C2 =>
                           REGISTERS_10_27_port, ZN => n15913);
   U14471 : OAI221_X1 port map( B1 => n10642, B2 => n13815, C1 => n10770, C2 =>
                           n303, A => n15914, ZN => n15909);
   U14472 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_27_port, B1 =>
                           n13819, B2 => REGISTERS_2_27_port, C1 => n360, C2 =>
                           REGISTERS_5_27_port, ZN => n15914);
   U14473 : OAI221_X1 port map( B1 => n10610, B2 => n13821, C1 => n11634, C2 =>
                           n304, A => n15915, ZN => n15908);
   U14474 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_27_port, B1 => 
                           n13825, B2 => REGISTERS_0_27_port, C1 => n13826, C2 
                           => REGISTERS_1_27_port, ZN => n15915);
   U14475 : NOR4_X1 port map( A1 => n15916, A2 => n15917, A3 => n15918, A4 => 
                           n15919, ZN => n15906);
   U14476 : OAI221_X1 port map( B1 => n11698, B2 => n362, C1 => n10962, C2 => 
                           n373, A => n15920, ZN => n15919);
   U14477 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_30_27_port, B1 => 
                           n395, B2 => REGISTERS_34_27_port, C1 => n406, C2 => 
                           REGISTERS_38_27_port, ZN => n15920);
   U14478 : OAI221_X1 port map( B1 => n11538, B2 => n417, C1 => n11666, C2 => 
                           n428, A => n15921, ZN => n15918);
   U14479 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_25_27_port, B1 => 
                           n450, B2 => REGISTERS_29_27_port, C1 => n461, C2 => 
                           REGISTERS_33_27_port, ZN => n15921);
   U14480 : OAI221_X1 port map( B1 => n11378, B2 => n472, C1 => n11506, C2 => 
                           n483, A => n15922, ZN => n15917);
   U14481 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_20_27_port, B1 => 
                           n505, B2 => REGISTERS_24_27_port, C1 => n516, C2 => 
                           REGISTERS_28_27_port, ZN => n15922);
   U14482 : OAI221_X1 port map( B1 => n11218, B2 => n527, C1 => n11346, C2 => 
                           n538, A => n15923, ZN => n15916);
   U14483 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_23_27_port, B1 => 
                           n560, B2 => REGISTERS_21_27_port, C1 => n571, C2 => 
                           REGISTERS_19_27_port, ZN => n15923);
   U14484 : NOR4_X1 port map( A1 => n15926, A2 => n15927, A3 => n15928, A4 => 
                           n15929, ZN => n15925);
   U14485 : OAI221_X1 port map( B1 => n11122, B2 => n307, C1 => n11058, C2 => 
                           n318, A => n15930, ZN => n15929);
   U14486 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_16_27_port, B1 => 
                           n119, B2 => REGISTERS_14_27_port, C1 => n13807, C2 
                           => REGISTERS_12_27_port, ZN => n15930);
   U14487 : OAI221_X1 port map( B1 => n11090, B2 => n13863, C1 => n10834, C2 =>
                           n13809, A => n15931, ZN => n15928);
   U14488 : AOI222_X1 port map( A1 => n340, A2 => REGISTERS_11_27_port, B1 => 
                           n13865, B2 => REGISTERS_9_27_port, C1 => n13813, C2 
                           => REGISTERS_7_27_port, ZN => n15931);
   U14489 : OAI221_X1 port map( B1 => n10930, B2 => n13866, C1 => n10674, C2 =>
                           n13815, A => n15932, ZN => n15927);
   U14490 : AOI222_X1 port map( A1 => n351, A2 => REGISTERS_6_27_port, B1 => 
                           n13868, B2 => REGISTERS_36_27_port, C1 => n13819, C2
                           => REGISTERS_3_27_port, ZN => n15932);
   U14491 : OAI221_X1 port map( B1 => n10770, B2 => n13869, C1 => n10642, C2 =>
                           n13821, A => n15933, ZN => n15926);
   U14492 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_27_port, B1 => 
                           n13871, B2 => REGISTERS_0_27_port, C1 => n13825, C2 
                           => REGISTERS_1_27_port, ZN => n15933);
   U14493 : NOR4_X1 port map( A1 => n15934, A2 => n15935, A3 => n15936, A4 => 
                           n15937, ZN => n15924);
   U14494 : OAI221_X1 port map( B1 => n11730, B2 => n362, C1 => n10994, C2 => 
                           n373, A => n15938, ZN => n15937);
   U14495 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_31_27_port, B1 => 
                           n395, B2 => REGISTERS_35_27_port, C1 => n406, C2 => 
                           REGISTERS_39_27_port, ZN => n15938);
   U14496 : OAI221_X1 port map( B1 => n11570, B2 => n417, C1 => n11698, C2 => 
                           n428, A => n15939, ZN => n15936);
   U14497 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_26_27_port, B1 => 
                           n450, B2 => REGISTERS_30_27_port, C1 => n461, C2 => 
                           REGISTERS_34_27_port, ZN => n15939);
   U14498 : OAI221_X1 port map( B1 => n11410, B2 => n472, C1 => n11538, C2 => 
                           n483, A => n15940, ZN => n15935);
   U14499 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_21_27_port, B1 => 
                           n505, B2 => REGISTERS_25_27_port, C1 => n516, C2 => 
                           REGISTERS_29_27_port, ZN => n15940);
   U14500 : OAI221_X1 port map( B1 => n11250, B2 => n527, C1 => n11378, C2 => 
                           n538, A => n15941, ZN => n15934);
   U14501 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_24_27_port, B1 => 
                           n560, B2 => REGISTERS_22_27_port, C1 => n571, C2 => 
                           REGISTERS_20_27_port, ZN => n15941);
   U14502 : AOI22_X1 port map( A1 => n13880, A2 => n5144, B1 => n13881, B2 => 
                           n5145, ZN => n15902);
   U14503 : NOR4_X1 port map( A1 => n15944, A2 => n15945, A3 => n15946, A4 => 
                           n15947, ZN => n15943);
   U14504 : OAI221_X1 port map( B1 => n11058, B2 => n307, C1 => n10994, C2 => 
                           n318, A => n15948, ZN => n15947);
   U14505 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_14_27_port, B1 => 
                           n13808, B2 => REGISTERS_38_27_port, C1 => n13889, C2
                           => REGISTERS_39_27_port, ZN => n15948);
   U14506 : OAI221_X1 port map( B1 => n10898, B2 => n13810, C1 => n10834, C2 =>
                           n13890, A => n15949, ZN => n15946);
   U14507 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_27_port, B1 => 
                           n346, B2 => REGISTERS_9_27_port, C1 => n13812, C2 =>
                           REGISTERS_16_27_port, ZN => n15949);
   U14508 : OAI221_X1 port map( B1 => n10738, B2 => n303, C1 => n10674, C2 => 
                           n13893, A => n15950, ZN => n15945);
   U14509 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_27_port, B1 => 
                           n357, B2 => REGISTERS_4_27_port, C1 => n13818, C2 =>
                           REGISTERS_11_27_port, ZN => n15950);
   U14510 : OAI221_X1 port map( B1 => n11602, B2 => n304, C1 => n10546, C2 => 
                           n13896, A => n15951, ZN => n15944);
   U14511 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_27_port, B1 => 
                           n13826, B2 => REGISTERS_0_27_port, C1 => n13824, C2 
                           => REGISTERS_6_27_port, ZN => n15951);
   U14512 : NOR4_X1 port map( A1 => n15952, A2 => n15953, A3 => n15954, A4 => 
                           n15955, ZN => n15942);
   U14513 : OAI221_X1 port map( B1 => n11666, B2 => n362, C1 => n10930, C2 => 
                           n373, A => n15956, ZN => n15955);
   U14514 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_29_27_port, B1 => 
                           n395, B2 => REGISTERS_33_27_port, C1 => n406, C2 => 
                           REGISTERS_37_27_port, ZN => n15956);
   U14515 : OAI221_X1 port map( B1 => n11506, B2 => n417, C1 => n11634, C2 => 
                           n428, A => n15957, ZN => n15954);
   U14516 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_24_27_port, B1 => 
                           n450, B2 => REGISTERS_28_27_port, C1 => n461, C2 => 
                           REGISTERS_32_27_port, ZN => n15957);
   U14517 : OAI221_X1 port map( B1 => n11346, B2 => n472, C1 => n11474, C2 => 
                           n483, A => n15958, ZN => n15953);
   U14518 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_19_27_port, B1 => 
                           n505, B2 => REGISTERS_23_27_port, C1 => n516, C2 => 
                           REGISTERS_27_27_port, ZN => n15958);
   U14519 : OAI221_X1 port map( B1 => n11186, B2 => n527, C1 => n11314, C2 => 
                           n538, A => n15959, ZN => n15952);
   U14520 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_22_27_port, B1 => 
                           n560, B2 => REGISTERS_20_27_port, C1 => n571, C2 => 
                           REGISTERS_18_27_port, ZN => n15959);
   U14521 : NOR4_X1 port map( A1 => n15962, A2 => n15963, A3 => n15964, A4 => 
                           n15965, ZN => n15961);
   U14522 : OAI221_X1 port map( B1 => n11026, B2 => n307, C1 => n10962, C2 => 
                           n318, A => n15966, ZN => n15965);
   U14523 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_13_27_port, B1 => 
                           n13808, B2 => REGISTERS_37_27_port, C1 => n13889, C2
                           => REGISTERS_38_27_port, ZN => n15966);
   U14524 : OAI221_X1 port map( B1 => n10866, B2 => n13810, C1 => n10802, C2 =>
                           n13890, A => n15967, ZN => n15964);
   U14525 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_27_port, B1 => 
                           n346, B2 => REGISTERS_8_27_port, C1 => n13812, C2 =>
                           REGISTERS_15_27_port, ZN => n15967);
   U14526 : OAI221_X1 port map( B1 => n10706, B2 => n303, C1 => n10642, C2 => 
                           n13893, A => n15968, ZN => n15963);
   U14527 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_27_port, B1 => 
                           n357, B2 => REGISTERS_3_27_port, C1 => n13818, C2 =>
                           REGISTERS_10_27_port, ZN => n15968);
   U14528 : OAI221_X1 port map( B1 => n11570, B2 => n304, C1 => n10460, C2 => 
                           n13896, A => n15969, ZN => n15962);
   U14529 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_27_port, B1 => 
                           n13917, B2 => REGISTERS_39_27_port, C1 => n13824, C2
                           => REGISTERS_5_27_port, ZN => n15969);
   U14530 : NOR4_X1 port map( A1 => n15970, A2 => n15971, A3 => n15972, A4 => 
                           n15973, ZN => n15960);
   U14531 : OAI221_X1 port map( B1 => n11634, B2 => n362, C1 => n10898, C2 => 
                           n373, A => n15974, ZN => n15973);
   U14532 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_28_27_port, B1 => 
                           n395, B2 => REGISTERS_32_27_port, C1 => n406, C2 => 
                           REGISTERS_36_27_port, ZN => n15974);
   U14533 : OAI221_X1 port map( B1 => n11474, B2 => n417, C1 => n11602, C2 => 
                           n428, A => n15975, ZN => n15972);
   U14534 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_23_27_port, B1 => 
                           n450, B2 => REGISTERS_27_27_port, C1 => n461, C2 => 
                           REGISTERS_31_27_port, ZN => n15975);
   U14535 : OAI221_X1 port map( B1 => n11314, B2 => n472, C1 => n11442, C2 => 
                           n483, A => n15976, ZN => n15971);
   U14536 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_18_27_port, B1 => 
                           n505, B2 => REGISTERS_22_27_port, C1 => n516, C2 => 
                           REGISTERS_26_27_port, ZN => n15976);
   U14537 : OAI221_X1 port map( B1 => n11154, B2 => n527, C1 => n11282, C2 => 
                           n538, A => n15977, ZN => n15970);
   U14538 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_21_27_port, B1 => 
                           n560, B2 => REGISTERS_19_27_port, C1 => n571, C2 => 
                           REGISTERS_17_27_port, ZN => n15977);
   U14539 : NAND3_X1 port map( A1 => n15978, A2 => n15979, A3 => n15980, ZN => 
                           n11876);
   U14540 : AOI221_X1 port map( B1 => n13792, B2 => n5149, C1 => n13793, C2 => 
                           MEM_IN(28), A => n15981, ZN => n15980);
   U14541 : OAI22_X1 port map( A1 => n10457, A2 => n251, B1 => n5151, B2 => 
                           n121, ZN => n15981);
   U14542 : NOR2_X1 port map( A1 => n5732, A2 => n13796, ZN => n5730);
   U14543 : INV_X1 port map( A => MEM_IN(28), ZN => n5732);
   U14544 : AOI22_X1 port map( A1 => n197, A2 => n5152, B1 => n150, B2 => n5153
                           , ZN => n15979);
   U14545 : NOR4_X1 port map( A1 => n15984, A2 => n15985, A3 => n15986, A4 => 
                           n15987, ZN => n15983);
   U14546 : OAI221_X1 port map( B1 => n11089, B2 => n307, C1 => n11025, C2 => 
                           n318, A => n15988, ZN => n15987);
   U14547 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_15_28_port, B1 => 
                           n13807, B2 => REGISTERS_11_28_port, C1 => n13808, C2
                           => REGISTERS_39_28_port, ZN => n15988);
   U14548 : OAI221_X1 port map( B1 => n10801, B2 => n13809, C1 => n10929, C2 =>
                           n13810, A => n15989, ZN => n15986);
   U14549 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_28_port, B1 =>
                           n13813, B2 => REGISTERS_6_28_port, C1 => n349, C2 =>
                           REGISTERS_10_28_port, ZN => n15989);
   U14550 : OAI221_X1 port map( B1 => n10641, B2 => n13815, C1 => n10769, C2 =>
                           n303, A => n15990, ZN => n15985);
   U14551 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_28_port, B1 =>
                           n13819, B2 => REGISTERS_2_28_port, C1 => n360, C2 =>
                           REGISTERS_5_28_port, ZN => n15990);
   U14552 : OAI221_X1 port map( B1 => n10609, B2 => n13821, C1 => n11633, C2 =>
                           n304, A => n15991, ZN => n15984);
   U14553 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_28_port, B1 => 
                           n13825, B2 => REGISTERS_0_28_port, C1 => n13826, C2 
                           => REGISTERS_1_28_port, ZN => n15991);
   U14554 : NOR4_X1 port map( A1 => n15992, A2 => n15993, A3 => n15994, A4 => 
                           n15995, ZN => n15982);
   U14555 : OAI221_X1 port map( B1 => n11697, B2 => n362, C1 => n10961, C2 => 
                           n373, A => n15996, ZN => n15995);
   U14556 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_30_28_port, B1 => 
                           n395, B2 => REGISTERS_34_28_port, C1 => n406, C2 => 
                           REGISTERS_38_28_port, ZN => n15996);
   U14557 : OAI221_X1 port map( B1 => n11537, B2 => n417, C1 => n11665, C2 => 
                           n428, A => n15997, ZN => n15994);
   U14558 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_25_28_port, B1 => 
                           n450, B2 => REGISTERS_29_28_port, C1 => n461, C2 => 
                           REGISTERS_33_28_port, ZN => n15997);
   U14559 : OAI221_X1 port map( B1 => n11377, B2 => n472, C1 => n11505, C2 => 
                           n483, A => n15998, ZN => n15993);
   U14560 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_20_28_port, B1 => 
                           n505, B2 => REGISTERS_24_28_port, C1 => n516, C2 => 
                           REGISTERS_28_28_port, ZN => n15998);
   U14561 : OAI221_X1 port map( B1 => n11217, B2 => n527, C1 => n11345, C2 => 
                           n538, A => n15999, ZN => n15992);
   U14562 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_23_28_port, B1 => 
                           n560, B2 => REGISTERS_21_28_port, C1 => n571, C2 => 
                           REGISTERS_19_28_port, ZN => n15999);
   U14563 : NOR4_X1 port map( A1 => n16002, A2 => n16003, A3 => n16004, A4 => 
                           n16005, ZN => n16001);
   U14564 : OAI221_X1 port map( B1 => n11121, B2 => n307, C1 => n11057, C2 => 
                           n318, A => n16006, ZN => n16005);
   U14565 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_16_28_port, B1 => 
                           n119, B2 => REGISTERS_14_28_port, C1 => n13807, C2 
                           => REGISTERS_12_28_port, ZN => n16006);
   U14566 : OAI221_X1 port map( B1 => n11089, B2 => n13863, C1 => n10833, C2 =>
                           n13809, A => n16007, ZN => n16004);
   U14567 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_28_port, B1 => 
                           n13865, B2 => REGISTERS_9_28_port, C1 => n13813, C2 
                           => REGISTERS_7_28_port, ZN => n16007);
   U14568 : OAI221_X1 port map( B1 => n10929, B2 => n13866, C1 => n10673, C2 =>
                           n13815, A => n16008, ZN => n16003);
   U14569 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_28_port, B1 => 
                           n13868, B2 => REGISTERS_36_28_port, C1 => n13819, C2
                           => REGISTERS_3_28_port, ZN => n16008);
   U14570 : OAI221_X1 port map( B1 => n10769, B2 => n13869, C1 => n10641, C2 =>
                           n13821, A => n16009, ZN => n16002);
   U14571 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_28_port, B1 => 
                           n13871, B2 => REGISTERS_0_28_port, C1 => n13825, C2 
                           => REGISTERS_1_28_port, ZN => n16009);
   U14572 : NOR4_X1 port map( A1 => n16010, A2 => n16011, A3 => n16012, A4 => 
                           n16013, ZN => n16000);
   U14573 : OAI221_X1 port map( B1 => n11729, B2 => n362, C1 => n10993, C2 => 
                           n373, A => n16014, ZN => n16013);
   U14574 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_31_28_port, B1 => 
                           n395, B2 => REGISTERS_35_28_port, C1 => n406, C2 => 
                           REGISTERS_39_28_port, ZN => n16014);
   U14575 : OAI221_X1 port map( B1 => n11569, B2 => n417, C1 => n11697, C2 => 
                           n428, A => n16015, ZN => n16012);
   U14576 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_26_28_port, B1 => 
                           n450, B2 => REGISTERS_30_28_port, C1 => n461, C2 => 
                           REGISTERS_34_28_port, ZN => n16015);
   U14577 : OAI221_X1 port map( B1 => n11409, B2 => n472, C1 => n11537, C2 => 
                           n483, A => n16016, ZN => n16011);
   U14578 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_21_28_port, B1 => 
                           n505, B2 => REGISTERS_25_28_port, C1 => n516, C2 => 
                           REGISTERS_29_28_port, ZN => n16016);
   U14579 : OAI221_X1 port map( B1 => n11249, B2 => n527, C1 => n11377, C2 => 
                           n538, A => n16017, ZN => n16010);
   U14580 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_24_28_port, B1 => 
                           n560, B2 => REGISTERS_22_28_port, C1 => n571, C2 => 
                           REGISTERS_20_28_port, ZN => n16017);
   U14581 : AOI22_X1 port map( A1 => n13880, A2 => n5154, B1 => n13881, B2 => 
                           n5155, ZN => n15978);
   U14582 : NOR4_X1 port map( A1 => n16020, A2 => n16021, A3 => n16022, A4 => 
                           n16023, ZN => n16019);
   U14583 : OAI221_X1 port map( B1 => n11057, B2 => n307, C1 => n10993, C2 => 
                           n318, A => n16024, ZN => n16023);
   U14584 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_14_28_port, B1 => 
                           n13808, B2 => REGISTERS_38_28_port, C1 => n13889, C2
                           => REGISTERS_39_28_port, ZN => n16024);
   U14585 : OAI221_X1 port map( B1 => n10897, B2 => n13810, C1 => n10833, C2 =>
                           n13890, A => n16025, ZN => n16022);
   U14586 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_28_port, B1 => 
                           n346, B2 => REGISTERS_9_28_port, C1 => n13812, C2 =>
                           REGISTERS_16_28_port, ZN => n16025);
   U14587 : OAI221_X1 port map( B1 => n10737, B2 => n303, C1 => n10673, C2 => 
                           n13893, A => n16026, ZN => n16021);
   U14588 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_28_port, B1 => 
                           n357, B2 => REGISTERS_4_28_port, C1 => n13818, C2 =>
                           REGISTERS_11_28_port, ZN => n16026);
   U14589 : OAI221_X1 port map( B1 => n11601, B2 => n304, C1 => n10545, C2 => 
                           n13896, A => n16027, ZN => n16020);
   U14590 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_28_port, B1 => 
                           n13826, B2 => REGISTERS_0_28_port, C1 => n13824, C2 
                           => REGISTERS_6_28_port, ZN => n16027);
   U14591 : NOR4_X1 port map( A1 => n16028, A2 => n16029, A3 => n16030, A4 => 
                           n16031, ZN => n16018);
   U14592 : OAI221_X1 port map( B1 => n11665, B2 => n362, C1 => n10929, C2 => 
                           n373, A => n16032, ZN => n16031);
   U14593 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_29_28_port, B1 => 
                           n395, B2 => REGISTERS_33_28_port, C1 => n406, C2 => 
                           REGISTERS_37_28_port, ZN => n16032);
   U14594 : OAI221_X1 port map( B1 => n11505, B2 => n417, C1 => n11633, C2 => 
                           n428, A => n16033, ZN => n16030);
   U14595 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_24_28_port, B1 => 
                           n450, B2 => REGISTERS_28_28_port, C1 => n461, C2 => 
                           REGISTERS_32_28_port, ZN => n16033);
   U14596 : OAI221_X1 port map( B1 => n11345, B2 => n472, C1 => n11473, C2 => 
                           n483, A => n16034, ZN => n16029);
   U14597 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_19_28_port, B1 => 
                           n505, B2 => REGISTERS_23_28_port, C1 => n516, C2 => 
                           REGISTERS_27_28_port, ZN => n16034);
   U14598 : OAI221_X1 port map( B1 => n11185, B2 => n527, C1 => n11313, C2 => 
                           n538, A => n16035, ZN => n16028);
   U14599 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_22_28_port, B1 => 
                           n560, B2 => REGISTERS_20_28_port, C1 => n571, C2 => 
                           REGISTERS_18_28_port, ZN => n16035);
   U14600 : NOR4_X1 port map( A1 => n16038, A2 => n16039, A3 => n16040, A4 => 
                           n16041, ZN => n16037);
   U14601 : OAI221_X1 port map( B1 => n11025, B2 => n307, C1 => n10961, C2 => 
                           n318, A => n16042, ZN => n16041);
   U14602 : AOI222_X1 port map( A1 => n329, A2 => REGISTERS_13_28_port, B1 => 
                           n13808, B2 => REGISTERS_37_28_port, C1 => n13889, C2
                           => REGISTERS_38_28_port, ZN => n16042);
   U14603 : OAI221_X1 port map( B1 => n10865, B2 => n13810, C1 => n10801, C2 =>
                           n13890, A => n16043, ZN => n16040);
   U14604 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_28_port, B1 => 
                           n346, B2 => REGISTERS_8_28_port, C1 => n13812, C2 =>
                           REGISTERS_15_28_port, ZN => n16043);
   U14605 : OAI221_X1 port map( B1 => n10705, B2 => n303, C1 => n10641, C2 => 
                           n13893, A => n16044, ZN => n16039);
   U14606 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_28_port, B1 => 
                           n357, B2 => REGISTERS_3_28_port, C1 => n13818, C2 =>
                           REGISTERS_10_28_port, ZN => n16044);
   U14607 : OAI221_X1 port map( B1 => n11569, B2 => n304, C1 => n10457, C2 => 
                           n13896, A => n16045, ZN => n16038);
   U14608 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_28_port, B1 => 
                           n13917, B2 => REGISTERS_39_28_port, C1 => n13824, C2
                           => REGISTERS_5_28_port, ZN => n16045);
   U14609 : NOR4_X1 port map( A1 => n16046, A2 => n16047, A3 => n16048, A4 => 
                           n16049, ZN => n16036);
   U14610 : OAI221_X1 port map( B1 => n11633, B2 => n362, C1 => n10897, C2 => 
                           n373, A => n16050, ZN => n16049);
   U14611 : AOI222_X1 port map( A1 => n384, A2 => REGISTERS_28_28_port, B1 => 
                           n395, B2 => REGISTERS_32_28_port, C1 => n406, C2 => 
                           REGISTERS_36_28_port, ZN => n16050);
   U14612 : OAI221_X1 port map( B1 => n11473, B2 => n417, C1 => n11601, C2 => 
                           n428, A => n16051, ZN => n16048);
   U14613 : AOI222_X1 port map( A1 => n439, A2 => REGISTERS_23_28_port, B1 => 
                           n450, B2 => REGISTERS_27_28_port, C1 => n461, C2 => 
                           REGISTERS_31_28_port, ZN => n16051);
   U14614 : OAI221_X1 port map( B1 => n11313, B2 => n472, C1 => n11441, C2 => 
                           n483, A => n16052, ZN => n16047);
   U14615 : AOI222_X1 port map( A1 => n494, A2 => REGISTERS_18_28_port, B1 => 
                           n505, B2 => REGISTERS_22_28_port, C1 => n516, C2 => 
                           REGISTERS_26_28_port, ZN => n16052);
   U14616 : OAI221_X1 port map( B1 => n11153, B2 => n527, C1 => n11281, C2 => 
                           n538, A => n16053, ZN => n16046);
   U14617 : AOI222_X1 port map( A1 => n549, A2 => REGISTERS_21_28_port, B1 => 
                           n560, B2 => REGISTERS_19_28_port, C1 => n571, C2 => 
                           REGISTERS_17_28_port, ZN => n16053);
   U14618 : NAND3_X1 port map( A1 => n16054, A2 => n16055, A3 => n16056, ZN => 
                           n11875);
   U14619 : AOI221_X1 port map( B1 => n13792, B2 => n5159, C1 => n13793, C2 => 
                           MEM_IN(29), A => n16057, ZN => n16056);
   U14620 : OAI22_X1 port map( A1 => n10454, A2 => n251, B1 => n5161, B2 => 
                           n121, ZN => n16057);
   U14621 : NOR2_X1 port map( A1 => n5739, A2 => n13796, ZN => n5737);
   U14622 : INV_X1 port map( A => MEM_IN(29), ZN => n5739);
   U14623 : AOI22_X1 port map( A1 => n197, A2 => n5162, B1 => n150, B2 => n5163
                           , ZN => n16055);
   U14624 : NOR4_X1 port map( A1 => n16060, A2 => n16061, A3 => n16062, A4 => 
                           n16063, ZN => n16059);
   U14625 : OAI221_X1 port map( B1 => n11088, B2 => n306, C1 => n11024, C2 => 
                           n317, A => n16064, ZN => n16063);
   U14626 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_15_29_port, B1 => 
                           n13807, B2 => REGISTERS_11_29_port, C1 => n13808, C2
                           => REGISTERS_39_29_port, ZN => n16064);
   U14627 : OAI221_X1 port map( B1 => n10800, B2 => n13809, C1 => n10928, C2 =>
                           n13810, A => n16065, ZN => n16062);
   U14628 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_29_port, B1 =>
                           n13813, B2 => REGISTERS_6_29_port, C1 => n349, C2 =>
                           REGISTERS_10_29_port, ZN => n16065);
   U14629 : OAI221_X1 port map( B1 => n10640, B2 => n13815, C1 => n10768, C2 =>
                           n303, A => n16066, ZN => n16061);
   U14630 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_29_port, B1 =>
                           n13819, B2 => REGISTERS_2_29_port, C1 => n360, C2 =>
                           REGISTERS_5_29_port, ZN => n16066);
   U14631 : OAI221_X1 port map( B1 => n10608, B2 => n13821, C1 => n11632, C2 =>
                           n304, A => n16067, ZN => n16060);
   U14632 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_29_port, B1 => 
                           n13825, B2 => REGISTERS_0_29_port, C1 => n13826, C2 
                           => REGISTERS_1_29_port, ZN => n16067);
   U14633 : NOR4_X1 port map( A1 => n16068, A2 => n16069, A3 => n16070, A4 => 
                           n16071, ZN => n16058);
   U14634 : OAI221_X1 port map( B1 => n11696, B2 => n361, C1 => n10960, C2 => 
                           n373, A => n16072, ZN => n16071);
   U14635 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_30_29_port, B1 => 
                           n394, B2 => REGISTERS_34_29_port, C1 => n405, C2 => 
                           REGISTERS_38_29_port, ZN => n16072);
   U14636 : OAI221_X1 port map( B1 => n11536, B2 => n416, C1 => n11664, C2 => 
                           n427, A => n16073, ZN => n16070);
   U14637 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_25_29_port, B1 => 
                           n449, B2 => REGISTERS_29_29_port, C1 => n460, C2 => 
                           REGISTERS_33_29_port, ZN => n16073);
   U14638 : OAI221_X1 port map( B1 => n11376, B2 => n471, C1 => n11504, C2 => 
                           n482, A => n16074, ZN => n16069);
   U14639 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_20_29_port, B1 => 
                           n504, B2 => REGISTERS_24_29_port, C1 => n515, C2 => 
                           REGISTERS_28_29_port, ZN => n16074);
   U14640 : OAI221_X1 port map( B1 => n11216, B2 => n526, C1 => n11344, C2 => 
                           n537, A => n16075, ZN => n16068);
   U14641 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_23_29_port, B1 => 
                           n559, B2 => REGISTERS_21_29_port, C1 => n570, C2 => 
                           REGISTERS_19_29_port, ZN => n16075);
   U14642 : NOR4_X1 port map( A1 => n16078, A2 => n16079, A3 => n16080, A4 => 
                           n16081, ZN => n16077);
   U14643 : OAI221_X1 port map( B1 => n11120, B2 => n306, C1 => n11056, C2 => 
                           n317, A => n16082, ZN => n16081);
   U14644 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_16_29_port, B1 => 
                           n119, B2 => REGISTERS_14_29_port, C1 => n13807, C2 
                           => REGISTERS_12_29_port, ZN => n16082);
   U14645 : OAI221_X1 port map( B1 => n11088, B2 => n13863, C1 => n10832, C2 =>
                           n13809, A => n16083, ZN => n16080);
   U14646 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_29_port, B1 => 
                           n13865, B2 => REGISTERS_9_29_port, C1 => n13813, C2 
                           => REGISTERS_7_29_port, ZN => n16083);
   U14647 : OAI221_X1 port map( B1 => n10928, B2 => n13866, C1 => n10672, C2 =>
                           n13815, A => n16084, ZN => n16079);
   U14648 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_29_port, B1 => 
                           n13868, B2 => REGISTERS_36_29_port, C1 => n13819, C2
                           => REGISTERS_3_29_port, ZN => n16084);
   U14649 : OAI221_X1 port map( B1 => n10768, B2 => n13869, C1 => n10640, C2 =>
                           n13821, A => n16085, ZN => n16078);
   U14650 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_29_port, B1 => 
                           n13871, B2 => REGISTERS_0_29_port, C1 => n13825, C2 
                           => REGISTERS_1_29_port, ZN => n16085);
   U14651 : NOR4_X1 port map( A1 => n16086, A2 => n16087, A3 => n16088, A4 => 
                           n16089, ZN => n16076);
   U14652 : OAI221_X1 port map( B1 => n11728, B2 => n361, C1 => n10992, C2 => 
                           n372, A => n16090, ZN => n16089);
   U14653 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_31_29_port, B1 => 
                           n394, B2 => REGISTERS_35_29_port, C1 => n405, C2 => 
                           REGISTERS_39_29_port, ZN => n16090);
   U14654 : OAI221_X1 port map( B1 => n11568, B2 => n416, C1 => n11696, C2 => 
                           n427, A => n16091, ZN => n16088);
   U14655 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_26_29_port, B1 => 
                           n449, B2 => REGISTERS_30_29_port, C1 => n460, C2 => 
                           REGISTERS_34_29_port, ZN => n16091);
   U14656 : OAI221_X1 port map( B1 => n11408, B2 => n471, C1 => n11536, C2 => 
                           n482, A => n16092, ZN => n16087);
   U14657 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_21_29_port, B1 => 
                           n504, B2 => REGISTERS_25_29_port, C1 => n515, C2 => 
                           REGISTERS_29_29_port, ZN => n16092);
   U14658 : OAI221_X1 port map( B1 => n11248, B2 => n526, C1 => n11376, C2 => 
                           n537, A => n16093, ZN => n16086);
   U14659 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_24_29_port, B1 => 
                           n559, B2 => REGISTERS_22_29_port, C1 => n570, C2 => 
                           REGISTERS_20_29_port, ZN => n16093);
   U14660 : AOI22_X1 port map( A1 => n13880, A2 => n5164, B1 => n13881, B2 => 
                           n5165, ZN => n16054);
   U14661 : NOR4_X1 port map( A1 => n16096, A2 => n16097, A3 => n16098, A4 => 
                           n16099, ZN => n16095);
   U14662 : OAI221_X1 port map( B1 => n11056, B2 => n306, C1 => n10992, C2 => 
                           n317, A => n16100, ZN => n16099);
   U14663 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_14_29_port, B1 => 
                           n13808, B2 => REGISTERS_38_29_port, C1 => n13889, C2
                           => REGISTERS_39_29_port, ZN => n16100);
   U14664 : OAI221_X1 port map( B1 => n10896, B2 => n13810, C1 => n10832, C2 =>
                           n13890, A => n16101, ZN => n16098);
   U14665 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_29_port, B1 => 
                           n346, B2 => REGISTERS_9_29_port, C1 => n13812, C2 =>
                           REGISTERS_16_29_port, ZN => n16101);
   U14666 : OAI221_X1 port map( B1 => n10736, B2 => n303, C1 => n10672, C2 => 
                           n13893, A => n16102, ZN => n16097);
   U14667 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_29_port, B1 => 
                           n357, B2 => REGISTERS_4_29_port, C1 => n13818, C2 =>
                           REGISTERS_11_29_port, ZN => n16102);
   U14668 : OAI221_X1 port map( B1 => n11600, B2 => n304, C1 => n10544, C2 => 
                           n13896, A => n16103, ZN => n16096);
   U14669 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_29_port, B1 => 
                           n13826, B2 => REGISTERS_0_29_port, C1 => n13824, C2 
                           => REGISTERS_6_29_port, ZN => n16103);
   U14670 : NOR4_X1 port map( A1 => n16104, A2 => n16105, A3 => n16106, A4 => 
                           n16107, ZN => n16094);
   U14671 : OAI221_X1 port map( B1 => n11664, B2 => n361, C1 => n10928, C2 => 
                           n372, A => n16108, ZN => n16107);
   U14672 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_29_29_port, B1 => 
                           n394, B2 => REGISTERS_33_29_port, C1 => n405, C2 => 
                           REGISTERS_37_29_port, ZN => n16108);
   U14673 : OAI221_X1 port map( B1 => n11504, B2 => n416, C1 => n11632, C2 => 
                           n427, A => n16109, ZN => n16106);
   U14674 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_24_29_port, B1 => 
                           n449, B2 => REGISTERS_28_29_port, C1 => n460, C2 => 
                           REGISTERS_32_29_port, ZN => n16109);
   U14675 : OAI221_X1 port map( B1 => n11344, B2 => n471, C1 => n11472, C2 => 
                           n482, A => n16110, ZN => n16105);
   U14676 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_19_29_port, B1 => 
                           n504, B2 => REGISTERS_23_29_port, C1 => n515, C2 => 
                           REGISTERS_27_29_port, ZN => n16110);
   U14677 : OAI221_X1 port map( B1 => n11184, B2 => n526, C1 => n11312, C2 => 
                           n537, A => n16111, ZN => n16104);
   U14678 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_22_29_port, B1 => 
                           n559, B2 => REGISTERS_20_29_port, C1 => n570, C2 => 
                           REGISTERS_18_29_port, ZN => n16111);
   U14679 : NOR4_X1 port map( A1 => n16114, A2 => n16115, A3 => n16116, A4 => 
                           n16117, ZN => n16113);
   U14680 : OAI221_X1 port map( B1 => n11024, B2 => n306, C1 => n10960, C2 => 
                           n317, A => n16118, ZN => n16117);
   U14681 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_13_29_port, B1 => 
                           n13808, B2 => REGISTERS_37_29_port, C1 => n13889, C2
                           => REGISTERS_38_29_port, ZN => n16118);
   U14682 : OAI221_X1 port map( B1 => n10864, B2 => n13810, C1 => n10800, C2 =>
                           n13890, A => n16119, ZN => n16116);
   U14683 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_29_port, B1 => 
                           n346, B2 => REGISTERS_8_29_port, C1 => n13812, C2 =>
                           REGISTERS_15_29_port, ZN => n16119);
   U14684 : OAI221_X1 port map( B1 => n10704, B2 => n303, C1 => n10640, C2 => 
                           n13893, A => n16120, ZN => n16115);
   U14685 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_29_port, B1 => 
                           n357, B2 => REGISTERS_3_29_port, C1 => n13818, C2 =>
                           REGISTERS_10_29_port, ZN => n16120);
   U14686 : OAI221_X1 port map( B1 => n11568, B2 => n304, C1 => n10454, C2 => 
                           n13896, A => n16121, ZN => n16114);
   U14687 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_29_port, B1 => 
                           n13917, B2 => REGISTERS_39_29_port, C1 => n13824, C2
                           => REGISTERS_5_29_port, ZN => n16121);
   U14688 : NOR4_X1 port map( A1 => n16122, A2 => n16123, A3 => n16124, A4 => 
                           n16125, ZN => n16112);
   U14689 : OAI221_X1 port map( B1 => n11632, B2 => n361, C1 => n10896, C2 => 
                           n372, A => n16126, ZN => n16125);
   U14690 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_28_29_port, B1 => 
                           n394, B2 => REGISTERS_32_29_port, C1 => n405, C2 => 
                           REGISTERS_36_29_port, ZN => n16126);
   U14691 : OAI221_X1 port map( B1 => n11472, B2 => n416, C1 => n11600, C2 => 
                           n427, A => n16127, ZN => n16124);
   U14692 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_23_29_port, B1 => 
                           n449, B2 => REGISTERS_27_29_port, C1 => n460, C2 => 
                           REGISTERS_31_29_port, ZN => n16127);
   U14693 : OAI221_X1 port map( B1 => n11312, B2 => n471, C1 => n11440, C2 => 
                           n482, A => n16128, ZN => n16123);
   U14694 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_18_29_port, B1 => 
                           n504, B2 => REGISTERS_22_29_port, C1 => n515, C2 => 
                           REGISTERS_26_29_port, ZN => n16128);
   U14695 : OAI221_X1 port map( B1 => n11152, B2 => n526, C1 => n11280, C2 => 
                           n537, A => n16129, ZN => n16122);
   U14696 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_21_29_port, B1 => 
                           n559, B2 => REGISTERS_19_29_port, C1 => n570, C2 => 
                           REGISTERS_17_29_port, ZN => n16129);
   U14697 : NAND3_X1 port map( A1 => n16130, A2 => n16131, A3 => n16132, ZN => 
                           n11874);
   U14698 : AOI221_X1 port map( B1 => n13792, B2 => n5169, C1 => n13793, C2 => 
                           MEM_IN(30), A => n16133, ZN => n16132);
   U14699 : OAI22_X1 port map( A1 => n10451, A2 => n251, B1 => n5171, B2 => 
                           n121, ZN => n16133);
   U14700 : NOR2_X1 port map( A1 => n5746, A2 => n13796, ZN => n5744);
   U14701 : INV_X1 port map( A => MEM_IN(30), ZN => n5746);
   U14702 : AOI22_X1 port map( A1 => n197, A2 => n5172, B1 => n150, B2 => n5173
                           , ZN => n16131);
   U14703 : NOR4_X1 port map( A1 => n16136, A2 => n16137, A3 => n16138, A4 => 
                           n16139, ZN => n16135);
   U14704 : OAI221_X1 port map( B1 => n11087, B2 => n306, C1 => n11023, C2 => 
                           n317, A => n16140, ZN => n16139);
   U14705 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_15_30_port, B1 => 
                           n13807, B2 => REGISTERS_11_30_port, C1 => n13808, C2
                           => REGISTERS_39_30_port, ZN => n16140);
   U14706 : OAI221_X1 port map( B1 => n10799, B2 => n13809, C1 => n10927, C2 =>
                           n13810, A => n16141, ZN => n16138);
   U14707 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_30_port, B1 =>
                           n13813, B2 => REGISTERS_6_30_port, C1 => n349, C2 =>
                           REGISTERS_10_30_port, ZN => n16141);
   U14708 : OAI221_X1 port map( B1 => n10639, B2 => n13815, C1 => n10767, C2 =>
                           n303, A => n16142, ZN => n16137);
   U14709 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_30_port, B1 =>
                           n13819, B2 => REGISTERS_2_30_port, C1 => n360, C2 =>
                           REGISTERS_5_30_port, ZN => n16142);
   U14710 : OAI221_X1 port map( B1 => n10607, B2 => n13821, C1 => n11631, C2 =>
                           n304, A => n16143, ZN => n16136);
   U14711 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_30_port, B1 => 
                           n13825, B2 => REGISTERS_0_30_port, C1 => n13826, C2 
                           => REGISTERS_1_30_port, ZN => n16143);
   U14712 : NOR4_X1 port map( A1 => n16144, A2 => n16145, A3 => n16146, A4 => 
                           n16147, ZN => n16134);
   U14713 : OAI221_X1 port map( B1 => n11695, B2 => n361, C1 => n10959, C2 => 
                           n372, A => n16148, ZN => n16147);
   U14714 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_30_30_port, B1 => 
                           n394, B2 => REGISTERS_34_30_port, C1 => n405, C2 => 
                           REGISTERS_38_30_port, ZN => n16148);
   U14715 : OAI221_X1 port map( B1 => n11535, B2 => n416, C1 => n11663, C2 => 
                           n427, A => n16149, ZN => n16146);
   U14716 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_25_30_port, B1 => 
                           n449, B2 => REGISTERS_29_30_port, C1 => n460, C2 => 
                           REGISTERS_33_30_port, ZN => n16149);
   U14717 : OAI221_X1 port map( B1 => n11375, B2 => n471, C1 => n11503, C2 => 
                           n482, A => n16150, ZN => n16145);
   U14718 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_20_30_port, B1 => 
                           n504, B2 => REGISTERS_24_30_port, C1 => n515, C2 => 
                           REGISTERS_28_30_port, ZN => n16150);
   U14719 : OAI221_X1 port map( B1 => n11215, B2 => n526, C1 => n11343, C2 => 
                           n537, A => n16151, ZN => n16144);
   U14720 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_23_30_port, B1 => 
                           n559, B2 => REGISTERS_21_30_port, C1 => n570, C2 => 
                           REGISTERS_19_30_port, ZN => n16151);
   U14721 : NOR4_X1 port map( A1 => n16154, A2 => n16155, A3 => n16156, A4 => 
                           n16157, ZN => n16153);
   U14722 : OAI221_X1 port map( B1 => n11119, B2 => n306, C1 => n11055, C2 => 
                           n317, A => n16158, ZN => n16157);
   U14723 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_16_30_port, B1 => 
                           n119, B2 => REGISTERS_14_30_port, C1 => n13807, C2 
                           => REGISTERS_12_30_port, ZN => n16158);
   U14724 : OAI221_X1 port map( B1 => n11087, B2 => n13863, C1 => n10831, C2 =>
                           n13809, A => n16159, ZN => n16156);
   U14725 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_30_port, B1 => 
                           n13865, B2 => REGISTERS_9_30_port, C1 => n13813, C2 
                           => REGISTERS_7_30_port, ZN => n16159);
   U14726 : OAI221_X1 port map( B1 => n10927, B2 => n13866, C1 => n10671, C2 =>
                           n13815, A => n16160, ZN => n16155);
   U14727 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_30_port, B1 => 
                           n13868, B2 => REGISTERS_36_30_port, C1 => n13819, C2
                           => REGISTERS_3_30_port, ZN => n16160);
   U14728 : OAI221_X1 port map( B1 => n10767, B2 => n13869, C1 => n10639, C2 =>
                           n13821, A => n16161, ZN => n16154);
   U14729 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_30_port, B1 => 
                           n13871, B2 => REGISTERS_0_30_port, C1 => n13825, C2 
                           => REGISTERS_1_30_port, ZN => n16161);
   U14730 : NOR4_X1 port map( A1 => n16162, A2 => n16163, A3 => n16164, A4 => 
                           n16165, ZN => n16152);
   U14731 : OAI221_X1 port map( B1 => n11727, B2 => n361, C1 => n10991, C2 => 
                           n372, A => n16166, ZN => n16165);
   U14732 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_31_30_port, B1 => 
                           n394, B2 => REGISTERS_35_30_port, C1 => n405, C2 => 
                           REGISTERS_39_30_port, ZN => n16166);
   U14733 : OAI221_X1 port map( B1 => n11567, B2 => n416, C1 => n11695, C2 => 
                           n427, A => n16167, ZN => n16164);
   U14734 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_26_30_port, B1 => 
                           n449, B2 => REGISTERS_30_30_port, C1 => n460, C2 => 
                           REGISTERS_34_30_port, ZN => n16167);
   U14735 : OAI221_X1 port map( B1 => n11407, B2 => n471, C1 => n11535, C2 => 
                           n482, A => n16168, ZN => n16163);
   U14736 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_21_30_port, B1 => 
                           n504, B2 => REGISTERS_25_30_port, C1 => n515, C2 => 
                           REGISTERS_29_30_port, ZN => n16168);
   U14737 : OAI221_X1 port map( B1 => n11247, B2 => n526, C1 => n11375, C2 => 
                           n537, A => n16169, ZN => n16162);
   U14738 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_24_30_port, B1 => 
                           n559, B2 => REGISTERS_22_30_port, C1 => n570, C2 => 
                           REGISTERS_20_30_port, ZN => n16169);
   U14739 : AOI22_X1 port map( A1 => n13880, A2 => n5174, B1 => n13881, B2 => 
                           n5175, ZN => n16130);
   U14740 : NOR4_X1 port map( A1 => n16172, A2 => n16173, A3 => n16174, A4 => 
                           n16175, ZN => n16171);
   U14741 : OAI221_X1 port map( B1 => n11055, B2 => n306, C1 => n10991, C2 => 
                           n317, A => n16176, ZN => n16175);
   U14742 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_14_30_port, B1 => 
                           n13808, B2 => REGISTERS_38_30_port, C1 => n13889, C2
                           => REGISTERS_39_30_port, ZN => n16176);
   U14743 : OAI221_X1 port map( B1 => n10895, B2 => n13810, C1 => n10831, C2 =>
                           n13890, A => n16177, ZN => n16174);
   U14744 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_30_port, B1 => 
                           n346, B2 => REGISTERS_9_30_port, C1 => n13812, C2 =>
                           REGISTERS_16_30_port, ZN => n16177);
   U14745 : OAI221_X1 port map( B1 => n10735, B2 => n303, C1 => n10671, C2 => 
                           n13893, A => n16178, ZN => n16173);
   U14746 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_30_port, B1 => 
                           n357, B2 => REGISTERS_4_30_port, C1 => n13818, C2 =>
                           REGISTERS_11_30_port, ZN => n16178);
   U14747 : OAI221_X1 port map( B1 => n11599, B2 => n304, C1 => n10543, C2 => 
                           n13896, A => n16179, ZN => n16172);
   U14748 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_30_port, B1 => 
                           n13826, B2 => REGISTERS_0_30_port, C1 => n13824, C2 
                           => REGISTERS_6_30_port, ZN => n16179);
   U14749 : NOR4_X1 port map( A1 => n16180, A2 => n16181, A3 => n16182, A4 => 
                           n16183, ZN => n16170);
   U14750 : OAI221_X1 port map( B1 => n11663, B2 => n361, C1 => n10927, C2 => 
                           n372, A => n16184, ZN => n16183);
   U14751 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_29_30_port, B1 => 
                           n394, B2 => REGISTERS_33_30_port, C1 => n405, C2 => 
                           REGISTERS_37_30_port, ZN => n16184);
   U14752 : OAI221_X1 port map( B1 => n11503, B2 => n416, C1 => n11631, C2 => 
                           n427, A => n16185, ZN => n16182);
   U14753 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_24_30_port, B1 => 
                           n449, B2 => REGISTERS_28_30_port, C1 => n460, C2 => 
                           REGISTERS_32_30_port, ZN => n16185);
   U14754 : OAI221_X1 port map( B1 => n11343, B2 => n471, C1 => n11471, C2 => 
                           n482, A => n16186, ZN => n16181);
   U14755 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_19_30_port, B1 => 
                           n504, B2 => REGISTERS_23_30_port, C1 => n515, C2 => 
                           REGISTERS_27_30_port, ZN => n16186);
   U14756 : OAI221_X1 port map( B1 => n11183, B2 => n526, C1 => n11311, C2 => 
                           n537, A => n16187, ZN => n16180);
   U14757 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_22_30_port, B1 => 
                           n559, B2 => REGISTERS_20_30_port, C1 => n570, C2 => 
                           REGISTERS_18_30_port, ZN => n16187);
   U14758 : NOR4_X1 port map( A1 => n16190, A2 => n16191, A3 => n16192, A4 => 
                           n16193, ZN => n16189);
   U14759 : OAI221_X1 port map( B1 => n11023, B2 => n306, C1 => n10959, C2 => 
                           n317, A => n16194, ZN => n16193);
   U14760 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_13_30_port, B1 => 
                           n13808, B2 => REGISTERS_37_30_port, C1 => n13889, C2
                           => REGISTERS_38_30_port, ZN => n16194);
   U14761 : OAI221_X1 port map( B1 => n10863, B2 => n13810, C1 => n10799, C2 =>
                           n13890, A => n16195, ZN => n16192);
   U14762 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_30_port, B1 => 
                           n346, B2 => REGISTERS_8_30_port, C1 => n13812, C2 =>
                           REGISTERS_15_30_port, ZN => n16195);
   U14763 : OAI221_X1 port map( B1 => n10703, B2 => n303, C1 => n10639, C2 => 
                           n13893, A => n16196, ZN => n16191);
   U14764 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_30_port, B1 => 
                           n357, B2 => REGISTERS_3_30_port, C1 => n13818, C2 =>
                           REGISTERS_10_30_port, ZN => n16196);
   U14765 : OAI221_X1 port map( B1 => n11567, B2 => n304, C1 => n10451, C2 => 
                           n13896, A => n16197, ZN => n16190);
   U14766 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_30_port, B1 => 
                           n13917, B2 => REGISTERS_39_30_port, C1 => n13824, C2
                           => REGISTERS_5_30_port, ZN => n16197);
   U14767 : NOR4_X1 port map( A1 => n16198, A2 => n16199, A3 => n16200, A4 => 
                           n16201, ZN => n16188);
   U14768 : OAI221_X1 port map( B1 => n11631, B2 => n361, C1 => n10895, C2 => 
                           n372, A => n16202, ZN => n16201);
   U14769 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_28_30_port, B1 => 
                           n394, B2 => REGISTERS_32_30_port, C1 => n405, C2 => 
                           REGISTERS_36_30_port, ZN => n16202);
   U14770 : OAI221_X1 port map( B1 => n11471, B2 => n416, C1 => n11599, C2 => 
                           n427, A => n16203, ZN => n16200);
   U14771 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_23_30_port, B1 => 
                           n449, B2 => REGISTERS_27_30_port, C1 => n460, C2 => 
                           REGISTERS_31_30_port, ZN => n16203);
   U14772 : OAI221_X1 port map( B1 => n11311, B2 => n471, C1 => n11439, C2 => 
                           n482, A => n16204, ZN => n16199);
   U14773 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_18_30_port, B1 => 
                           n504, B2 => REGISTERS_22_30_port, C1 => n515, C2 => 
                           REGISTERS_26_30_port, ZN => n16204);
   U14774 : OAI221_X1 port map( B1 => n11151, B2 => n526, C1 => n11279, C2 => 
                           n537, A => n16205, ZN => n16198);
   U14775 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_21_30_port, B1 => 
                           n559, B2 => REGISTERS_19_30_port, C1 => n570, C2 => 
                           REGISTERS_17_30_port, ZN => n16205);
   U14776 : NAND3_X1 port map( A1 => n16206, A2 => n16207, A3 => n16208, ZN => 
                           n11873);
   U14777 : AOI221_X1 port map( B1 => n13792, B2 => n5179, C1 => n13793, C2 => 
                           MEM_IN(31), A => n16209, ZN => n16208);
   U14778 : OAI22_X1 port map( A1 => n10448, A2 => n251, B1 => n5181, B2 => 
                           n121, ZN => n16209);
   U14779 : NOR2_X1 port map( A1 => n5753, A2 => n13796, ZN => n5751);
   U14780 : INV_X1 port map( A => MEM_IN(31), ZN => n5753);
   U14781 : NAND2_X1 port map( A1 => n5206, A2 => n13632, ZN => n13628);
   U14782 : NAND2_X1 port map( A1 => n13337, A2 => n5206, ZN => n13632);
   U14783 : AOI22_X1 port map( A1 => n197, A2 => n5191, B1 => n150, B2 => n5192
                           , ZN => n16207);
   U14784 : NOR4_X1 port map( A1 => n16216, A2 => n16217, A3 => n16218, A4 => 
                           n16219, ZN => n16215);
   U14785 : OAI221_X1 port map( B1 => n11086, B2 => n306, C1 => n11022, C2 => 
                           n317, A => n16220, ZN => n16219);
   U14786 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_15_31_port, B1 => 
                           n13807, B2 => REGISTERS_11_31_port, C1 => n13808, C2
                           => REGISTERS_39_31_port, ZN => n16220);
   U14787 : OAI221_X1 port map( B1 => n10798, B2 => n13809, C1 => n10926, C2 =>
                           n13810, A => n16221, ZN => n16218);
   U14788 : AOI222_X1 port map( A1 => n13812, A2 => REGISTERS_17_31_port, B1 =>
                           n13813, B2 => REGISTERS_6_31_port, C1 => n347, C2 =>
                           REGISTERS_10_31_port, ZN => n16221);
   U14789 : OAI221_X1 port map( B1 => n10638, B2 => n13815, C1 => n10766, C2 =>
                           n303, A => n16222, ZN => n16217);
   U14790 : AOI222_X1 port map( A1 => n13818, A2 => REGISTERS_12_31_port, B1 =>
                           n13819, B2 => REGISTERS_2_31_port, C1 => n358, C2 =>
                           REGISTERS_5_31_port, ZN => n16222);
   U14791 : OAI221_X1 port map( B1 => n10606, B2 => n13821, C1 => n11630, C2 =>
                           n304, A => n16223, ZN => n16216);
   U14792 : AOI222_X1 port map( A1 => n13824, A2 => REGISTERS_7_31_port, B1 => 
                           n13825, B2 => REGISTERS_0_31_port, C1 => n13826, C2 
                           => REGISTERS_1_31_port, ZN => n16223);
   U14793 : NOR4_X1 port map( A1 => n16224, A2 => n16225, A3 => n16226, A4 => 
                           n16227, ZN => n16214);
   U14794 : OAI221_X1 port map( B1 => n11694, B2 => n361, C1 => n10958, C2 => 
                           n372, A => n16228, ZN => n16227);
   U14795 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_30_31_port, B1 => 
                           n394, B2 => REGISTERS_34_31_port, C1 => n405, C2 => 
                           REGISTERS_38_31_port, ZN => n16228);
   U14796 : OAI221_X1 port map( B1 => n11534, B2 => n416, C1 => n11662, C2 => 
                           n427, A => n16229, ZN => n16226);
   U14797 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_25_31_port, B1 => 
                           n449, B2 => REGISTERS_29_31_port, C1 => n460, C2 => 
                           REGISTERS_33_31_port, ZN => n16229);
   U14798 : OAI221_X1 port map( B1 => n11374, B2 => n471, C1 => n11502, C2 => 
                           n482, A => n16230, ZN => n16225);
   U14799 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_20_31_port, B1 => 
                           n504, B2 => REGISTERS_24_31_port, C1 => n515, C2 => 
                           REGISTERS_28_31_port, ZN => n16230);
   U14800 : OAI221_X1 port map( B1 => n11214, B2 => n526, C1 => n11342, C2 => 
                           n537, A => n16231, ZN => n16224);
   U14801 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_23_31_port, B1 => 
                           n559, B2 => REGISTERS_21_31_port, C1 => n570, C2 => 
                           REGISTERS_19_31_port, ZN => n16231);
   U14802 : INV_X1 port map( A => n13787, ZN => n13781);
   U14803 : NOR2_X1 port map( A1 => n13485, A2 => n4787, ZN => n13787);
   U14804 : NOR4_X1 port map( A1 => n16235, A2 => n16236, A3 => n16237, A4 => 
                           n16238, ZN => n16234);
   U14805 : OAI221_X1 port map( B1 => n11118, B2 => n306, C1 => n11054, C2 => 
                           n317, A => n16239, ZN => n16238);
   U14806 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_16_31_port, B1 => 
                           n119, B2 => REGISTERS_14_31_port, C1 => n13807, C2 
                           => REGISTERS_12_31_port, ZN => n16239);
   U14807 : INV_X1 port map( A => n13810, ZN => n13862_port);
   U14808 : OAI221_X1 port map( B1 => n11086, B2 => n13863, C1 => n10830, C2 =>
                           n13809, A => n16240, ZN => n16237);
   U14809 : AOI222_X1 port map( A1 => n339, A2 => REGISTERS_11_31_port, B1 => 
                           n13865, B2 => REGISTERS_9_31_port, C1 => n13813, C2 
                           => REGISTERS_7_31_port, ZN => n16240);
   U14810 : OAI221_X1 port map( B1 => n10926, B2 => n13866, C1 => n10670, C2 =>
                           n13815, A => n16241, ZN => n16236);
   U14811 : AOI222_X1 port map( A1 => n350, A2 => REGISTERS_6_31_port, B1 => 
                           n13868, B2 => REGISTERS_36_31_port, C1 => n13819, C2
                           => REGISTERS_3_31_port, ZN => n16241);
   U14812 : OAI221_X1 port map( B1 => n10766, B2 => n13869, C1 => n10638, C2 =>
                           n13821, A => n16242, ZN => n16235);
   U14813 : AOI222_X1 port map( A1 => n13826, A2 => REGISTERS_2_31_port, B1 => 
                           n13871, B2 => REGISTERS_0_31_port, C1 => n13825, C2 
                           => REGISTERS_1_31_port, ZN => n16242);
   U14814 : NOR4_X1 port map( A1 => n16246, A2 => n16247, A3 => n16248, A4 => 
                           n16249, ZN => n16233);
   U14815 : OAI221_X1 port map( B1 => n11726, B2 => n361, C1 => n10990, C2 => 
                           n372, A => n16250, ZN => n16249);
   U14816 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_31_31_port, B1 => 
                           n394, B2 => REGISTERS_35_31_port, C1 => n405, C2 => 
                           REGISTERS_39_31_port, ZN => n16250);
   U14817 : OAI221_X1 port map( B1 => n11566, B2 => n416, C1 => n11694, C2 => 
                           n427, A => n16251, ZN => n16248);
   U14818 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_26_31_port, B1 => 
                           n449, B2 => REGISTERS_30_31_port, C1 => n460, C2 => 
                           REGISTERS_34_31_port, ZN => n16251);
   U14819 : OAI221_X1 port map( B1 => n11406, B2 => n471, C1 => n11534, C2 => 
                           n482, A => n16252, ZN => n16247);
   U14820 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_21_31_port, B1 => 
                           n504, B2 => REGISTERS_25_31_port, C1 => n515, C2 => 
                           REGISTERS_29_31_port, ZN => n16252);
   U14821 : OAI221_X1 port map( B1 => n11246, B2 => n526, C1 => n11374, C2 => 
                           n537, A => n16253, ZN => n16246);
   U14822 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_24_31_port, B1 => 
                           n559, B2 => REGISTERS_22_31_port, C1 => n570, C2 => 
                           REGISTERS_20_31_port, ZN => n16253);
   U14823 : OR2_X1 port map( A1 => n13490, A2 => n4787, ZN => n16213);
   U14824 : AOI22_X1 port map( A1 => n13880, A2 => n5195, B1 => n13881, B2 => 
                           n5196, ZN => n16206);
   U14825 : NOR4_X1 port map( A1 => n16256, A2 => n16257, A3 => n16258, A4 => 
                           n16259, ZN => n16255);
   U14826 : OAI221_X1 port map( B1 => n11054, B2 => n306, C1 => n10990, C2 => 
                           n317, A => n16260, ZN => n16259);
   U14827 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_14_31_port, B1 => 
                           n13808, B2 => REGISTERS_38_31_port, C1 => n13889, C2
                           => REGISTERS_39_31_port, ZN => n16260);
   U14828 : OAI221_X1 port map( B1 => n10894, B2 => n13810, C1 => n10830, C2 =>
                           n13890, A => n16261, ZN => n16258);
   U14829 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_8_31_port, B1 => 
                           n341, B2 => REGISTERS_9_31_port, C1 => n13812, C2 =>
                           REGISTERS_16_31_port, ZN => n16261);
   U14830 : OAI221_X1 port map( B1 => n10734, B2 => n303, C1 => n10670, C2 => 
                           n13893, A => n16262, ZN => n16257);
   U14831 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_3_31_port, B1 => 
                           n352, B2 => REGISTERS_4_31_port, C1 => n13818, C2 =>
                           REGISTERS_11_31_port, ZN => n16262);
   U14832 : OAI221_X1 port map( B1 => n11598, B2 => n304, C1 => n10542, C2 => 
                           n13896, A => n16263, ZN => n16256);
   U14833 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_2_31_port, B1 => 
                           n13826, B2 => REGISTERS_0_31_port, C1 => n13824, C2 
                           => REGISTERS_6_31_port, ZN => n16263);
   U14834 : NOR3_X1 port map( A1 => n11842, A2 => n11859, A3 => CWP_3_port, ZN 
                           => n16244);
   U14835 : NOR4_X1 port map( A1 => n16265, A2 => n16266, A3 => n16267, A4 => 
                           n16268, ZN => n16254);
   U14836 : OAI221_X1 port map( B1 => n11662, B2 => n361, C1 => n10926, C2 => 
                           n372, A => n16269, ZN => n16268);
   U14837 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_29_31_port, B1 => 
                           n394, B2 => REGISTERS_33_31_port, C1 => n405, C2 => 
                           REGISTERS_37_31_port, ZN => n16269);
   U14838 : OAI221_X1 port map( B1 => n11502, B2 => n416, C1 => n11630, C2 => 
                           n427, A => n16270, ZN => n16267);
   U14839 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_24_31_port, B1 => 
                           n449, B2 => REGISTERS_28_31_port, C1 => n460, C2 => 
                           REGISTERS_32_31_port, ZN => n16270);
   U14840 : OAI221_X1 port map( B1 => n11342, B2 => n471, C1 => n11470, C2 => 
                           n482, A => n16271, ZN => n16266);
   U14841 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_19_31_port, B1 => 
                           n504, B2 => REGISTERS_23_31_port, C1 => n515, C2 => 
                           REGISTERS_27_31_port, ZN => n16271);
   U14842 : OAI221_X1 port map( B1 => n11182, B2 => n526, C1 => n11310, C2 => 
                           n537, A => n16272, ZN => n16265);
   U14843 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_22_31_port, B1 => 
                           n559, B2 => REGISTERS_20_31_port, C1 => n570, C2 => 
                           REGISTERS_18_31_port, ZN => n16272);
   U14844 : NOR2_X1 port map( A1 => n11858, A2 => n4787, ZN => n13633);
   U14845 : NOR4_X1 port map( A1 => n16275, A2 => n16276, A3 => n16277, A4 => 
                           n16278, ZN => n16274);
   U14846 : OAI221_X1 port map( B1 => n11022, B2 => n306, C1 => n10958, C2 => 
                           n317, A => n16279, ZN => n16278);
   U14847 : AOI222_X1 port map( A1 => n328, A2 => REGISTERS_13_31_port, B1 => 
                           n13808, B2 => REGISTERS_37_31_port, C1 => n13889, C2
                           => REGISTERS_38_31_port, ZN => n16279);
   U14848 : AND2_X1 port map( A1 => n16245, A2 => n16281, ZN => n13806);
   U14849 : NAND2_X1 port map( A1 => n16243, A2 => n16281, ZN => n13804);
   U14850 : NAND2_X1 port map( A1 => n16282, A2 => n16283, ZN => n13803);
   U14851 : OAI221_X1 port map( B1 => n10862, B2 => n13810, C1 => n10798, C2 =>
                           n13890, A => n16284, ZN => n16277);
   U14852 : AOI222_X1 port map( A1 => n13892, A2 => REGISTERS_7_31_port, B1 => 
                           n344, B2 => REGISTERS_8_31_port, C1 => n13812, C2 =>
                           REGISTERS_15_31_port, ZN => n16284);
   U14853 : AND2_X1 port map( A1 => n16283, A2 => n16281, ZN => n13814);
   U14854 : OAI221_X1 port map( B1 => n10702, B2 => n303, C1 => n10638, C2 => 
                           n13893, A => n16288, ZN => n16276);
   U14855 : AOI222_X1 port map( A1 => n13895, A2 => REGISTERS_2_31_port, B1 => 
                           n355, B2 => REGISTERS_3_31_port, C1 => n13818, C2 =>
                           REGISTERS_10_31_port, ZN => n16288);
   U14856 : AND2_X1 port map( A1 => n16287, A2 => n16285, ZN => n13820);
   U14857 : OAI221_X1 port map( B1 => n11566, B2 => n304, C1 => n10448, C2 => 
                           n13896, A => n16291, ZN => n16275);
   U14858 : AOI222_X1 port map( A1 => n13898, A2 => REGISTERS_1_31_port, B1 => 
                           n13917, B2 => REGISTERS_39_31_port, C1 => n13824, C2
                           => REGISTERS_5_31_port, ZN => n16291);
   U14859 : AND2_X1 port map( A1 => n16292, A2 => CWP_5_port, ZN => n16285);
   U14860 : NOR4_X1 port map( A1 => n16293, A2 => n16294, A3 => n16295, A4 => 
                           n16296, ZN => n16273);
   U14861 : OAI221_X1 port map( B1 => n11630, B2 => n361, C1 => n10894, C2 => 
                           n372, A => n16297, ZN => n16296);
   U14862 : AOI222_X1 port map( A1 => n383, A2 => REGISTERS_28_31_port, B1 => 
                           n394, B2 => REGISTERS_32_31_port, C1 => n405, C2 => 
                           REGISTERS_36_31_port, ZN => n16297);
   U14863 : AND2_X1 port map( A1 => n16280, A2 => n16290, ZN => n13836_port);
   U14864 : AND2_X1 port map( A1 => n16283, A2 => n16280, ZN => n13835_port);
   U14865 : AND2_X1 port map( A1 => n16298, A2 => n16290, ZN => n13834_port);
   U14866 : NAND2_X1 port map( A1 => n16287, A2 => n16280, ZN => n13831_port);
   U14867 : OAI221_X1 port map( B1 => n11470, B2 => n416, C1 => n11598, C2 => 
                           n427, A => n16299, ZN => n16295);
   U14868 : AOI222_X1 port map( A1 => n438, A2 => REGISTERS_23_31_port, B1 => 
                           n449, B2 => REGISTERS_27_31_port, C1 => n460, C2 => 
                           REGISTERS_31_31_port, ZN => n16299);
   U14869 : AND2_X1 port map( A1 => n16298, A2 => n16264, ZN => n13842_port);
   U14870 : AND2_X1 port map( A1 => n16298, A2 => n16287, ZN => n13841_port);
   U14871 : AND2_X1 port map( A1 => n16282, A2 => n16264, ZN => n13840_port);
   U14872 : NOR2_X1 port map( A1 => n16300, A2 => n11862, ZN => n16264);
   U14873 : NAND2_X1 port map( A1 => n16289, A2 => n16280, ZN => n13838_port);
   U14874 : AND2_X1 port map( A1 => n11842, A2 => n16292, ZN => n16280);
   U14875 : NAND2_X1 port map( A1 => n16298, A2 => n16243, ZN => n13837_port);
   U14876 : OAI221_X1 port map( B1 => n11310, B2 => n471, C1 => n11438, C2 => 
                           n482, A => n16301, ZN => n16294);
   U14877 : AOI222_X1 port map( A1 => n493, A2 => REGISTERS_18_31_port, B1 => 
                           n504, B2 => REGISTERS_22_31_port, C1 => n515, C2 => 
                           REGISTERS_26_31_port, ZN => n16301);
   U14878 : AND2_X1 port map( A1 => n16298, A2 => n16289, ZN => n13848_port);
   U14879 : AND2_X1 port map( A1 => n16282, A2 => n16243, ZN => n13847_port);
   U14880 : NOR3_X1 port map( A1 => n11861, A2 => n11862, A3 => CWP_0_port, ZN 
                           => n16243);
   U14881 : AND2_X1 port map( A1 => n16282, A2 => n16289, ZN => n13846_port);
   U14882 : NOR3_X1 port map( A1 => CWP_0_port, A2 => n11862, A3 => CWP_2_port,
                           ZN => n16289);
   U14883 : NAND2_X1 port map( A1 => n16298, A2 => n16245, ZN => n13844_port);
   U14884 : NAND2_X1 port map( A1 => n16298, A2 => n16286, ZN => n13843_port);
   U14885 : OAI221_X1 port map( B1 => n11150, B2 => n526, C1 => n11278, C2 => 
                           n537, A => n16302, ZN => n16293);
   U14886 : AOI222_X1 port map( A1 => n548, A2 => REGISTERS_21_31_port, B1 => 
                           n559, B2 => REGISTERS_19_31_port, C1 => n570, C2 => 
                           REGISTERS_17_31_port, ZN => n16302);
   U14887 : AND2_X1 port map( A1 => n16282, A2 => n16286, ZN => n13854_port);
   U14888 : AND2_X1 port map( A1 => n16282, A2 => n16287, ZN => n13853_port);
   U14889 : NOR3_X1 port map( A1 => n11862, A2 => n11863, A3 => CWP_2_port, ZN 
                           => n16287);
   U14890 : AND2_X1 port map( A1 => n16282, A2 => n16245, ZN => n13852_port);
   U14891 : NOR2_X1 port map( A1 => n16300, A2 => CWP_1_port, ZN => n16245);
   U14892 : NAND2_X1 port map( A1 => n16298, A2 => n16283, ZN => n13850_port);
   U14893 : NOR3_X1 port map( A1 => CWP_0_port, A2 => CWP_1_port, A3 => 
                           CWP_2_port, ZN => n16283);
   U14894 : NOR3_X1 port map( A1 => CWP_5_port, A2 => n11859, A3 => CWP_3_port,
                           ZN => n16298);
   U14895 : NAND2_X1 port map( A1 => n16282, A2 => n16290, ZN => n13849_port);
   U14896 : NOR3_X1 port map( A1 => CWP_5_port, A2 => n11860, A3 => CWP_4_port,
                           ZN => n16282);
   U14897 : INV_X1 port map( A => n16232, ZN => n16212);
   U14898 : AOI22_X1 port map( A1 => n16303, A2 => n16210, B1 => n4841, B2 => 
                           n251, ZN => n16232);
   U14899 : INV_X1 port map( A => n208, ZN => n4841);
   U14900 : AND3_X1 port map( A1 => n208, A2 => n251, A3 => n16304, ZN => 
                           n16210);
   U14901 : OAI22_X1 port map( A1 => n4786, A2 => n16305, B1 => n16306, B2 => 
                           n5204, ZN => n13795);
   U14902 : INV_X1 port map( A => n4843, ZN => n4788);
   U14903 : NAND3_X1 port map( A1 => n4810, A2 => ENABLE, A3 => n300, ZN => 
                           n4843);
   U14904 : INV_X1 port map( A => n16307, ZN => n4810);
   U14905 : NOR2_X1 port map( A1 => n10078, A2 => n16211, ZN => n16306);
   U14906 : INV_X1 port map( A => n16303, ZN => n16211);
   U14907 : INV_X1 port map( A => n16304, ZN => n10078);
   U14908 : AOI21_X1 port map( B1 => n13642, B2 => n10226, A => n13638, ZN => 
                           n16304);
   U14909 : OR2_X1 port map( A1 => n5775, A2 => n5926, ZN => n13642);
   U14910 : NOR3_X1 port map( A1 => n11868, A2 => n11869, A3 => n1, ZN => n5926
                           );
   U14911 : AOI221_X1 port map( B1 => n10073, B2 => n7558, C1 => n5206, C2 => 
                           n13638, A => RESET, ZN => n16305);
   U14912 : NAND2_X1 port map( A1 => n11871, A2 => n13337, ZN => n13638);
   U14913 : AND2_X1 port map( A1 => n11858, A2 => n11855, ZN => n13337);
   U14914 : NAND2_X1 port map( A1 => n10226, A2 => n5215, ZN => n11858);
   U14915 : AND2_X1 port map( A1 => n13490, A2 => n13485, ZN => n11871);
   U14916 : NAND2_X1 port map( A1 => n10226, A2 => n5372, ZN => n13485);
   U14917 : NAND2_X1 port map( A1 => n10226, A2 => n5526, ZN => n13490);
   U14918 : INV_X1 port map( A => n6374, ZN => n7558);
   U14919 : NAND3_X1 port map( A1 => n10076, A2 => n10077, A3 => n10075, ZN => 
                           n6374);
   U14920 : INV_X1 port map( A => n11857, ZN => n10075);
   U14921 : INV_X1 port map( A => n10225, ZN => n10077);
   U14922 : INV_X1 port map( A => n13339, ZN => n10073);
   U14923 : NAND3_X1 port map( A1 => n8742, A2 => n8743, A3 => n7560, ZN => 
                           n13339);
   U14924 : AND2_X1 port map( A1 => WR, A2 => n6376, ZN => n7560);
   U14925 : AOI21_X1 port map( B1 => n5775, B2 => n16308, A => n13788, ZN => 
                           n16303);
   U14926 : OAI221_X1 port map( B1 => n13643, B2 => n13341, C1 => n16309, C2 =>
                           n16310, A => n13640, ZN => n13788);
   U14927 : AOI21_X1 port map( B1 => n5372, B2 => n16308, A => n16311, ZN => 
                           n13640);
   U14928 : INV_X1 port map( A => n13491, ZN => n16311);
   U14929 : AOI22_X1 port map( A1 => n6381, A2 => n10226, B1 => n5215, B2 => 
                           n16308, ZN => n13491);
   U14930 : NOR3_X1 port map( A1 => n11868, A2 => n11869, A3 => n11867, ZN => 
                           n5215);
   U14931 : NOR3_X1 port map( A1 => n11867, A2 => n11868, A3 => n808, ZN => 
                           n5372);
   U14932 : INV_X1 port map( A => n5526, ZN => n16309);
   U14933 : NOR3_X1 port map( A1 => n11867, A2 => n11869, A3 => n839, ZN => 
                           n5526);
   U14934 : INV_X1 port map( A => n10226, ZN => n13341);
   U14935 : NOR2_X1 port map( A1 => n6079, A2 => n6228, ZN => n13643);
   U14936 : NOR3_X1 port map( A1 => n840, A2 => n11869, A3 => n1, ZN => n6228);
   U14937 : NOR3_X1 port map( A1 => n807, A2 => n11868, A3 => n1, ZN => n6079);
   U14938 : INV_X1 port map( A => n16310, ZN => n16308);
   U14939 : NAND3_X1 port map( A1 => SWP_5_port, A2 => SWP_4_port, A3 => n11866
                           , ZN => n16310);
   U14940 : NOR2_X1 port map( A1 => n11855, A2 => n4787, ZN => n13482);
   U14941 : NAND2_X1 port map( A1 => n10080, A2 => n6381, ZN => n11855);
   U14942 : NOR3_X1 port map( A1 => n813, A2 => n814, A3 => n1, ZN => n6381);
   U14943 : MUX2_X1 port map( A => FILL_port, B => n16312, S => n16313, Z => 
                           n11872);
   U14944 : NOR2_X1 port map( A1 => n4786, A2 => n4846, ZN => n16313);
   U14945 : MUX2_X1 port map( A => n13796, B => n4847, S => n2, Z => n16312);
   U14946 : OAI21_X1 port map( B1 => CALL, B2 => n117, A => n16307, ZN => n4847
                           );
   U14947 : NAND4_X1 port map( A1 => n16315, A2 => n16316, A3 => n16317, A4 => 
                           n16318, ZN => n16307);
   U14948 : NOR4_X1 port map( A1 => n16319, A2 => CWP_30_port, A3 => 
                           CWP_29_port, A4 => CWP_28_port, ZN => n16318);
   U14949 : NOR4_X1 port map( A1 => CWP_27_port, A2 => CWP_26_port, A3 => 
                           CWP_25_port, A4 => CWP_24_port, ZN => n16317);
   U14950 : NOR4_X1 port map( A1 => CWP_23_port, A2 => CWP_22_port, A3 => 
                           CWP_9_port, A4 => CWP_8_port, ZN => n16316);
   U14951 : NOR4_X1 port map( A1 => CWP_7_port, A2 => CWP_6_port, A3 => 
                           CWP_31_port, A4 => n372, ZN => n16315);
   U14952 : NAND2_X1 port map( A1 => n16290, A2 => n16281, ZN => n13832_port);
   U14953 : NOR3_X1 port map( A1 => CWP_1_port, A2 => n11861, A3 => CWP_0_port,
                           ZN => n16290);
   U14954 : OAI21_X1 port map( B1 => n10413, B2 => n210, A => n16320, ZN => 
                           n11816);
   U14955 : AOI22_X1 port map( A1 => N50368, A2 => n207, B1 => N12268, B2 => 
                           n214, ZN => n16320);
   U14956 : OAI21_X1 port map( B1 => n10412, B2 => n210, A => n16321, ZN => 
                           n11815);
   U14957 : AOI22_X1 port map( A1 => N50367, A2 => n207, B1 => N12267, B2 => 
                           n214, ZN => n16321);
   U14958 : OAI21_X1 port map( B1 => n10411, B2 => n210, A => n16322, ZN => 
                           n11814);
   U14959 : AOI22_X1 port map( A1 => N50366, A2 => n207, B1 => N12266, B2 => 
                           n214, ZN => n16322);
   U14960 : OAI21_X1 port map( B1 => n10410, B2 => n210, A => n16323, ZN => 
                           n11813);
   U14961 : AOI22_X1 port map( A1 => N50365, A2 => n207, B1 => N12265, B2 => 
                           n214, ZN => n16323);
   U14962 : OAI21_X1 port map( B1 => n10409, B2 => n210, A => n16324, ZN => 
                           n11812);
   U14963 : AOI22_X1 port map( A1 => N50364, A2 => n207, B1 => N12264, B2 => 
                           n214, ZN => n16324);
   U14964 : OAI21_X1 port map( B1 => n10408, B2 => n210, A => n16325, ZN => 
                           n11811);
   U14965 : AOI22_X1 port map( A1 => N50363, A2 => n207, B1 => N12263, B2 => 
                           n214, ZN => n16325);
   U14966 : OAI21_X1 port map( B1 => n10407, B2 => n210, A => n16326, ZN => 
                           n11810);
   U14967 : AOI22_X1 port map( A1 => N50362, A2 => n207, B1 => N12262, B2 => 
                           n214, ZN => n16326);
   U14968 : OAI21_X1 port map( B1 => n10406, B2 => n210, A => n16327, ZN => 
                           n11809);
   U14969 : AOI22_X1 port map( A1 => N50361, A2 => n207, B1 => N12261, B2 => 
                           n214, ZN => n16327);
   U14970 : OAI21_X1 port map( B1 => n10405, B2 => n210, A => n16328, ZN => 
                           n11808);
   U14971 : AOI22_X1 port map( A1 => N50360, A2 => n207, B1 => N12260, B2 => 
                           n214, ZN => n16328);
   U14972 : OAI21_X1 port map( B1 => n10404, B2 => n210, A => n16329, ZN => 
                           n11807);
   U14973 : AOI22_X1 port map( A1 => N50359, A2 => n207, B1 => N12259, B2 => 
                           n214, ZN => n16329);
   U14974 : OAI21_X1 port map( B1 => n10403, B2 => n210, A => n16330, ZN => 
                           n11806);
   U14975 : AOI22_X1 port map( A1 => N50358, A2 => n207, B1 => N12258, B2 => 
                           n214, ZN => n16330);
   U14976 : OAI21_X1 port map( B1 => n10402, B2 => n210, A => n16331, ZN => 
                           n11805);
   U14977 : AOI22_X1 port map( A1 => N50357, A2 => n207, B1 => N12257, B2 => 
                           n214, ZN => n16331);
   U14978 : OAI21_X1 port map( B1 => n10401, B2 => n210, A => n16332, ZN => 
                           n11804);
   U14979 : AOI22_X1 port map( A1 => N50356, A2 => n207, B1 => N12256, B2 => 
                           n214, ZN => n16332);
   U14980 : OAI21_X1 port map( B1 => n10400, B2 => n210, A => n16333, ZN => 
                           n11803);
   U14981 : AOI22_X1 port map( A1 => N50355, A2 => n207, B1 => N12255, B2 => 
                           n214, ZN => n16333);
   U14982 : OAI21_X1 port map( B1 => n10399, B2 => n210, A => n16334, ZN => 
                           n11802);
   U14983 : AOI22_X1 port map( A1 => N50354, A2 => n207, B1 => N12254, B2 => 
                           n214, ZN => n16334);
   U14984 : OAI21_X1 port map( B1 => n10398, B2 => n210, A => n16335, ZN => 
                           n11801);
   U14985 : AOI22_X1 port map( A1 => N50353, A2 => n207, B1 => N12253, B2 => 
                           n214, ZN => n16335);
   U14986 : OAI21_X1 port map( B1 => n10397, B2 => n210, A => n16336, ZN => 
                           n11800);
   U14987 : AOI22_X1 port map( A1 => N50352, A2 => n207, B1 => N12252, B2 => 
                           n214, ZN => n16336);
   U14988 : OAI21_X1 port map( B1 => n10396, B2 => n210, A => n16337, ZN => 
                           n11799);
   U14989 : AOI22_X1 port map( A1 => N50351, A2 => n207, B1 => N12251, B2 => 
                           n214, ZN => n16337);
   U14990 : OAI21_X1 port map( B1 => n10395, B2 => n210, A => n16338, ZN => 
                           n11798);
   U14991 : AOI22_X1 port map( A1 => N50350, A2 => n207, B1 => N12250, B2 => 
                           n214, ZN => n16338);
   U14992 : OAI21_X1 port map( B1 => n10394, B2 => n210, A => n16339, ZN => 
                           n11797);
   U14993 : AOI22_X1 port map( A1 => N50349, A2 => n207, B1 => N12249, B2 => 
                           n214, ZN => n16339);
   U14994 : OAI21_X1 port map( B1 => n10393, B2 => n210, A => n16340, ZN => 
                           n11796);
   U14995 : AOI22_X1 port map( A1 => N50348, A2 => n207, B1 => N12248, B2 => 
                           n214, ZN => n16340);
   U14996 : OAI21_X1 port map( B1 => n10392, B2 => n210, A => n16341, ZN => 
                           n11795);
   U14997 : AOI22_X1 port map( A1 => N50347, A2 => n207, B1 => N12247, B2 => 
                           n214, ZN => n16341);
   U14998 : OAI21_X1 port map( B1 => n10391, B2 => n210, A => n16342, ZN => 
                           n11794);
   U14999 : AOI22_X1 port map( A1 => N50346, A2 => n207, B1 => N12246, B2 => 
                           n214, ZN => n16342);
   U15000 : OAI21_X1 port map( B1 => n10390, B2 => n210, A => n16343, ZN => 
                           n11793);
   U15001 : AOI22_X1 port map( A1 => N50345, A2 => n207, B1 => N12245, B2 => 
                           n214, ZN => n16343);
   U15002 : OAI21_X1 port map( B1 => n10389, B2 => n210, A => n16344, ZN => 
                           n11792);
   U15003 : AOI22_X1 port map( A1 => N50344, A2 => n207, B1 => N12244, B2 => 
                           n214, ZN => n16344);
   U15004 : OAI21_X1 port map( B1 => n10388, B2 => n210, A => n16345, ZN => 
                           n11791);
   U15005 : AOI22_X1 port map( A1 => N50343, A2 => n207, B1 => N12243, B2 => 
                           n214, ZN => n16345);
   U15006 : OAI21_X1 port map( B1 => n4786, B2 => n4809, A => n4752, ZN => 
                           n4851);
   U15007 : OAI21_X1 port map( B1 => n4844, B2 => n116, A => n4787, ZN => 
                           n16346);
   U15008 : INV_X1 port map( A => n4784, ZN => n4785);
   U15009 : NOR2_X1 port map( A1 => n4844, A2 => n16455, ZN => n4784);
   U15010 : OAI21_X1 port map( B1 => n16347, B2 => n16348, A => n11790, ZN => 
                           n4840);
   U15011 : NAND2_X1 port map( A1 => n16349, A2 => n16350, ZN => n16348);
   U15012 : NOR4_X1 port map( A1 => CWP_8_port, A2 => CWP_7_port, A3 => 
                           CWP_6_port, A4 => CWP_5_port, ZN => n16349);
   U15013 : NAND4_X1 port map( A1 => n11818, A2 => n11817, A3 => n16351, A4 => 
                           n16352, ZN => n16347);
   U15014 : AOI21_X1 port map( B1 => n16292, B2 => CWP_2_port, A => n16319, ZN 
                           => n16351);
   U15015 : NOR2_X1 port map( A1 => n11859, A2 => n11860, ZN => n16292);
   U15016 : INV_X1 port map( A => CALL, ZN => n4844);
   U15017 : INV_X1 port map( A => n4812, ZN => n4809);
   U15018 : NOR2_X1 port map( A1 => n16314, A2 => n2, ZN => n4812);
   U15019 : INV_X1 port map( A => RET, ZN => n4846);
   U15020 : NAND2_X1 port map( A1 => n11790, A2 => n16353, ZN => n16314);
   U15021 : NAND4_X1 port map( A1 => n16354, A2 => n16350, A3 => n16352, A4 => 
                           n16355, ZN => n16353);
   U15022 : NOR4_X1 port map( A1 => n16319, A2 => n16356, A3 => CWP_30_port, A4
                           => CWP_29_port, ZN => n16355);
   U15023 : OAI21_X1 port map( B1 => n11862, B2 => n11861, A => n16300, ZN => 
                           n16356);
   U15024 : NAND2_X1 port map( A1 => CWP_2_port, A2 => CWP_0_port, ZN => n16300
                           );
   U15025 : NAND4_X1 port map( A1 => n16357, A2 => n16358, A3 => n16359, A4 => 
                           n16360, ZN => n16319);
   U15026 : AND3_X1 port map( A1 => n11828, A2 => n11826, A3 => n11827, ZN => 
                           n16360);
   U15027 : AND3_X1 port map( A1 => n11831, A2 => n11829, A3 => n11830, ZN => 
                           n16359);
   U15028 : AND3_X1 port map( A1 => n11834, A2 => n11832, A3 => n11833, ZN => 
                           n16358);
   U15029 : AND3_X1 port map( A1 => n11837, A2 => n11835, A3 => n11836, ZN => 
                           n16357);
   U15030 : NOR4_X1 port map( A1 => CWP_28_port, A2 => CWP_27_port, A3 => 
                           CWP_26_port, A4 => CWP_25_port, ZN => n16352);
   U15031 : NOR4_X1 port map( A1 => CWP_24_port, A2 => CWP_23_port, A3 => 
                           CWP_22_port, A4 => CWP_9_port, ZN => n16350);
   U15032 : AND4_X1 port map( A1 => n11839, A2 => n11840, A3 => n11841, A4 => 
                           n16281, ZN => n16354);
   U15033 : OAI221_X1 port map( B1 => n5536, B2 => n16361, C1 => n10355, C2 => 
                           n16362, A => n16363, ZN => n10540);
   U15034 : NAND2_X1 port map( A1 => N4526, A2 => n16364, ZN => n16363);
   U15035 : OAI221_X1 port map( B1 => n5536, B2 => n16365, C1 => n10323, C2 => 
                           n16366, A => n16367, ZN => n10539);
   U15036 : NAND2_X1 port map( A1 => N4420, A2 => n16368, ZN => n16367);
   U15037 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n5368, ZN => n5536);
   U15038 : OAI221_X1 port map( B1 => n5544, B2 => n16361, C1 => n10356, C2 => 
                           n16362, A => n16369, ZN => n10537);
   U15039 : NAND2_X1 port map( A1 => N4525, A2 => n16364, ZN => n16369);
   U15040 : OAI221_X1 port map( B1 => n5544, B2 => n16365, C1 => n10324, C2 => 
                           n16366, A => n16370, ZN => n10536);
   U15041 : NAND2_X1 port map( A1 => N4419, A2 => n16368, ZN => n16370);
   U15042 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n5368, ZN => n5544);
   U15043 : OAI221_X1 port map( B1 => n5551, B2 => n16361, C1 => n10357, C2 => 
                           n16362, A => n16371, ZN => n10534);
   U15044 : NAND2_X1 port map( A1 => N4524, A2 => n16364, ZN => n16371);
   U15045 : OAI221_X1 port map( B1 => n5551, B2 => n16365, C1 => n10325, C2 => 
                           n16366, A => n16372, ZN => n10533);
   U15046 : NAND2_X1 port map( A1 => N4418, A2 => n16368, ZN => n16372);
   U15047 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n5368, ZN => n5551);
   U15048 : OAI221_X1 port map( B1 => n5558, B2 => n16361, C1 => n10358, C2 => 
                           n16362, A => n16373, ZN => n10531);
   U15049 : NAND2_X1 port map( A1 => N4523, A2 => n16364, ZN => n16373);
   U15050 : OAI221_X1 port map( B1 => n5558, B2 => n16365, C1 => n10326, C2 => 
                           n16366, A => n16374, ZN => n10530);
   U15051 : NAND2_X1 port map( A1 => N4417, A2 => n16368, ZN => n16374);
   U15052 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n5368, ZN => n5558);
   U15053 : OAI221_X1 port map( B1 => n5565, B2 => n16361, C1 => n10359, C2 => 
                           n16362, A => n16375, ZN => n10528);
   U15054 : NAND2_X1 port map( A1 => N4522, A2 => n16364, ZN => n16375);
   U15055 : OAI221_X1 port map( B1 => n5565, B2 => n16365, C1 => n10327, C2 => 
                           n16366, A => n16376, ZN => n10527);
   U15056 : NAND2_X1 port map( A1 => N4416, A2 => n16368, ZN => n16376);
   U15057 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n5368, ZN => n5565);
   U15058 : OAI221_X1 port map( B1 => n5572, B2 => n16361, C1 => n10360, C2 => 
                           n16362, A => n16377, ZN => n10525);
   U15059 : NAND2_X1 port map( A1 => N4521, A2 => n16364, ZN => n16377);
   U15060 : OAI221_X1 port map( B1 => n5572, B2 => n16365, C1 => n10328, C2 => 
                           n16366, A => n16378, ZN => n10524);
   U15061 : NAND2_X1 port map( A1 => N4415, A2 => n16368, ZN => n16378);
   U15062 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n5368, ZN => n5572);
   U15063 : OAI221_X1 port map( B1 => n5579, B2 => n16361, C1 => n10361, C2 => 
                           n16362, A => n16379, ZN => n10522);
   U15064 : NAND2_X1 port map( A1 => N4520, A2 => n16364, ZN => n16379);
   U15065 : OAI221_X1 port map( B1 => n5579, B2 => n16365, C1 => n10329, C2 => 
                           n16366, A => n16380, ZN => n10521);
   U15066 : NAND2_X1 port map( A1 => N4414, A2 => n16368, ZN => n16380);
   U15067 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n5368, ZN => n5579);
   U15068 : OAI221_X1 port map( B1 => n5586, B2 => n16361, C1 => n10362, C2 => 
                           n16362, A => n16381, ZN => n10519);
   U15069 : NAND2_X1 port map( A1 => N4519, A2 => n16364, ZN => n16381);
   U15070 : OAI221_X1 port map( B1 => n5586, B2 => n16365, C1 => n10330, C2 => 
                           n16366, A => n16382, ZN => n10518);
   U15071 : NAND2_X1 port map( A1 => N4413, A2 => n16368, ZN => n16382);
   U15072 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n5368, ZN => n5586);
   U15073 : OAI221_X1 port map( B1 => n5593, B2 => n16361, C1 => n10363, C2 => 
                           n16362, A => n16383, ZN => n10516);
   U15074 : NAND2_X1 port map( A1 => N4518, A2 => n16364, ZN => n16383);
   U15075 : OAI221_X1 port map( B1 => n5593, B2 => n16365, C1 => n10331, C2 => 
                           n16366, A => n16384, ZN => n10515);
   U15076 : NAND2_X1 port map( A1 => N4412, A2 => n16368, ZN => n16384);
   U15077 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n5368, ZN => n5593);
   U15078 : OAI221_X1 port map( B1 => n5600, B2 => n16361, C1 => n10364, C2 => 
                           n16362, A => n16385, ZN => n10513);
   U15079 : NAND2_X1 port map( A1 => N4517, A2 => n16364, ZN => n16385);
   U15080 : OAI221_X1 port map( B1 => n5600, B2 => n16365, C1 => n10332, C2 => 
                           n16366, A => n16386, ZN => n10512);
   U15081 : NAND2_X1 port map( A1 => N4411, A2 => n16368, ZN => n16386);
   U15082 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n5368, ZN => n5600);
   U15083 : OAI221_X1 port map( B1 => n5607, B2 => n16361, C1 => n10365, C2 => 
                           n16362, A => n16387, ZN => n10510);
   U15084 : NAND2_X1 port map( A1 => N4516, A2 => n16364, ZN => n16387);
   U15085 : OAI221_X1 port map( B1 => n5607, B2 => n16365, C1 => n10333, C2 => 
                           n16366, A => n16388, ZN => n10509);
   U15086 : NAND2_X1 port map( A1 => N4410, A2 => n16368, ZN => n16388);
   U15087 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n5368, ZN => n5607);
   U15088 : OAI221_X1 port map( B1 => n5614, B2 => n16361, C1 => n10366, C2 => 
                           n16362, A => n16389, ZN => n10507);
   U15089 : NAND2_X1 port map( A1 => N4515, A2 => n16364, ZN => n16389);
   U15090 : OAI221_X1 port map( B1 => n5614, B2 => n16365, C1 => n10334, C2 => 
                           n16366, A => n16390, ZN => n10506);
   U15091 : NAND2_X1 port map( A1 => N4409, A2 => n16368, ZN => n16390);
   U15092 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n5368, ZN => n5614);
   U15093 : OAI221_X1 port map( B1 => n5621, B2 => n16361, C1 => n10367, C2 => 
                           n16362, A => n16391, ZN => n10504);
   U15094 : NAND2_X1 port map( A1 => N4514, A2 => n16364, ZN => n16391);
   U15095 : OAI221_X1 port map( B1 => n5621, B2 => n16365, C1 => n10335, C2 => 
                           n16366, A => n16392, ZN => n10503);
   U15096 : NAND2_X1 port map( A1 => N4408, A2 => n16368, ZN => n16392);
   U15097 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n5368, ZN => n5621);
   U15098 : OAI221_X1 port map( B1 => n5628, B2 => n16361, C1 => n10368, C2 => 
                           n16362, A => n16393, ZN => n10501);
   U15099 : NAND2_X1 port map( A1 => N4513, A2 => n16364, ZN => n16393);
   U15100 : OAI221_X1 port map( B1 => n5628, B2 => n16365, C1 => n10336, C2 => 
                           n16366, A => n16394, ZN => n10500);
   U15101 : NAND2_X1 port map( A1 => N4407, A2 => n16368, ZN => n16394);
   U15102 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n5368, ZN => n5628);
   U15103 : OAI221_X1 port map( B1 => n5635, B2 => n16361, C1 => n10369, C2 => 
                           n16362, A => n16395, ZN => n10498);
   U15104 : NAND2_X1 port map( A1 => N4512, A2 => n16364, ZN => n16395);
   U15105 : OAI221_X1 port map( B1 => n5635, B2 => n16365, C1 => n10337, C2 => 
                           n16366, A => n16396, ZN => n10497);
   U15106 : NAND2_X1 port map( A1 => N4406, A2 => n16368, ZN => n16396);
   U15107 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n5368, ZN => n5635);
   U15108 : OAI221_X1 port map( B1 => n5642, B2 => n16361, C1 => n10370, C2 => 
                           n16362, A => n16397, ZN => n10495);
   U15109 : NAND2_X1 port map( A1 => N4511, A2 => n16364, ZN => n16397);
   U15110 : OAI221_X1 port map( B1 => n5642, B2 => n16365, C1 => n10338, C2 => 
                           n16366, A => n16398, ZN => n10494);
   U15111 : NAND2_X1 port map( A1 => N4405, A2 => n16368, ZN => n16398);
   U15112 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n5368, ZN => n5642);
   U15113 : OAI221_X1 port map( B1 => n5649, B2 => n16361, C1 => n10371, C2 => 
                           n16362, A => n16399, ZN => n10492);
   U15114 : NAND2_X1 port map( A1 => N4510, A2 => n16364, ZN => n16399);
   U15115 : OAI221_X1 port map( B1 => n5649, B2 => n16365, C1 => n10339, C2 => 
                           n16366, A => n16400, ZN => n10491);
   U15116 : NAND2_X1 port map( A1 => N4404, A2 => n16368, ZN => n16400);
   U15117 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n5368, ZN => n5649);
   U15118 : OAI221_X1 port map( B1 => n5656, B2 => n16361, C1 => n10372, C2 => 
                           n16362, A => n16401, ZN => n10489);
   U15119 : NAND2_X1 port map( A1 => N4509, A2 => n16364, ZN => n16401);
   U15120 : OAI221_X1 port map( B1 => n5656, B2 => n16365, C1 => n10340, C2 => 
                           n16366, A => n16402, ZN => n10488);
   U15121 : NAND2_X1 port map( A1 => N4403, A2 => n16368, ZN => n16402);
   U15122 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n5368, ZN => n5656);
   U15123 : OAI221_X1 port map( B1 => n5663, B2 => n16361, C1 => n10373, C2 => 
                           n16362, A => n16403, ZN => n10486);
   U15124 : NAND2_X1 port map( A1 => N4508, A2 => n16364, ZN => n16403);
   U15125 : OAI221_X1 port map( B1 => n5663, B2 => n16365, C1 => n10341, C2 => 
                           n16366, A => n16404, ZN => n10485);
   U15126 : NAND2_X1 port map( A1 => N4402, A2 => n16368, ZN => n16404);
   U15127 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n5368, ZN => n5663);
   U15128 : OAI221_X1 port map( B1 => n5670, B2 => n16361, C1 => n10374, C2 => 
                           n16362, A => n16405, ZN => n10483);
   U15129 : NAND2_X1 port map( A1 => N4507, A2 => n16364, ZN => n16405);
   U15130 : OAI221_X1 port map( B1 => n5670, B2 => n16365, C1 => n10342, C2 => 
                           n16366, A => n16406, ZN => n10482);
   U15131 : NAND2_X1 port map( A1 => N4401, A2 => n16368, ZN => n16406);
   U15132 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n5368, ZN => n5670);
   U15133 : OAI221_X1 port map( B1 => n5677, B2 => n16361, C1 => n10375, C2 => 
                           n16362, A => n16407, ZN => n10480);
   U15134 : NAND2_X1 port map( A1 => N4506, A2 => n16364, ZN => n16407);
   U15135 : OAI221_X1 port map( B1 => n5677, B2 => n16365, C1 => n10343, C2 => 
                           n16366, A => n16408, ZN => n10479);
   U15136 : NAND2_X1 port map( A1 => N4400, A2 => n16368, ZN => n16408);
   U15137 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n5368, ZN => n5677);
   U15138 : OAI221_X1 port map( B1 => n5684, B2 => n16361, C1 => n10376, C2 => 
                           n16362, A => n16409, ZN => n10477);
   U15139 : NAND2_X1 port map( A1 => N4505, A2 => n16364, ZN => n16409);
   U15140 : OAI221_X1 port map( B1 => n5684, B2 => n16365, C1 => n10344, C2 => 
                           n16366, A => n16410, ZN => n10476);
   U15141 : NAND2_X1 port map( A1 => N4399, A2 => n16368, ZN => n16410);
   U15142 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n5368, ZN => n5684);
   U15143 : OAI221_X1 port map( B1 => n5691, B2 => n16361, C1 => n10377, C2 => 
                           n16362, A => n16411, ZN => n10474);
   U15144 : NAND2_X1 port map( A1 => N4504, A2 => n16364, ZN => n16411);
   U15145 : OAI221_X1 port map( B1 => n5691, B2 => n16365, C1 => n10345, C2 => 
                           n16366, A => n16412, ZN => n10473);
   U15146 : NAND2_X1 port map( A1 => N4398, A2 => n16368, ZN => n16412);
   U15147 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n5368, ZN => n5691);
   U15148 : OAI221_X1 port map( B1 => n5698, B2 => n16361, C1 => n10378, C2 => 
                           n16362, A => n16413, ZN => n10471);
   U15149 : NAND2_X1 port map( A1 => N4503, A2 => n16364, ZN => n16413);
   U15150 : OAI221_X1 port map( B1 => n5698, B2 => n16365, C1 => n10346, C2 => 
                           n16366, A => n16414, ZN => n10470);
   U15151 : NAND2_X1 port map( A1 => N4397, A2 => n16368, ZN => n16414);
   U15152 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n5368, ZN => n5698);
   U15153 : OAI221_X1 port map( B1 => n5705, B2 => n16361, C1 => n10379, C2 => 
                           n16362, A => n16415, ZN => n10468);
   U15154 : NAND2_X1 port map( A1 => N4502, A2 => n16364, ZN => n16415);
   U15155 : OAI221_X1 port map( B1 => n5705, B2 => n16365, C1 => n10347, C2 => 
                           n16366, A => n16416, ZN => n10467);
   U15156 : NAND2_X1 port map( A1 => N4396, A2 => n16368, ZN => n16416);
   U15157 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n5368, ZN => n5705);
   U15158 : OAI221_X1 port map( B1 => n5712, B2 => n16361, C1 => n10380, C2 => 
                           n16362, A => n16417, ZN => n10465);
   U15159 : NAND2_X1 port map( A1 => N4501, A2 => n16364, ZN => n16417);
   U15160 : OAI221_X1 port map( B1 => n5712, B2 => n16365, C1 => n10348, C2 => 
                           n16366, A => n16418, ZN => n10464);
   U15161 : NAND2_X1 port map( A1 => N4395, A2 => n16368, ZN => n16418);
   U15162 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n5368, ZN => n5712);
   U15163 : OAI221_X1 port map( B1 => n5719, B2 => n16361, C1 => n10381, C2 => 
                           n16362, A => n16419, ZN => n10462);
   U15164 : NAND2_X1 port map( A1 => N4500, A2 => n16364, ZN => n16419);
   U15165 : OAI221_X1 port map( B1 => n5719, B2 => n16365, C1 => n10349, C2 => 
                           n16366, A => n16420, ZN => n10461);
   U15166 : NAND2_X1 port map( A1 => N4394, A2 => n16368, ZN => n16420);
   U15167 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n5368, ZN => n5719);
   U15168 : OAI221_X1 port map( B1 => n5726, B2 => n16361, C1 => n10382, C2 => 
                           n16362, A => n16421, ZN => n10459);
   U15169 : NAND2_X1 port map( A1 => N4499, A2 => n16364, ZN => n16421);
   U15170 : OAI221_X1 port map( B1 => n5726, B2 => n16365, C1 => n10350, C2 => 
                           n16366, A => n16422, ZN => n10458);
   U15171 : NAND2_X1 port map( A1 => N4393, A2 => n16368, ZN => n16422);
   U15172 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n5368, ZN => n5726);
   U15173 : OAI221_X1 port map( B1 => n5733, B2 => n16361, C1 => n10383, C2 => 
                           n16362, A => n16423, ZN => n10456);
   U15174 : NAND2_X1 port map( A1 => N4498, A2 => n16364, ZN => n16423);
   U15175 : OAI221_X1 port map( B1 => n5733, B2 => n16365, C1 => n10351, C2 => 
                           n16366, A => n16424, ZN => n10455);
   U15176 : NAND2_X1 port map( A1 => N4392, A2 => n16368, ZN => n16424);
   U15177 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n5368, ZN => n5733);
   U15178 : OAI221_X1 port map( B1 => n5740, B2 => n16361, C1 => n10384, C2 => 
                           n16362, A => n16425, ZN => n10453);
   U15179 : NAND2_X1 port map( A1 => N4497, A2 => n16364, ZN => n16425);
   U15180 : OAI221_X1 port map( B1 => n5740, B2 => n16365, C1 => n10352, C2 => 
                           n16366, A => n16426, ZN => n10452);
   U15181 : NAND2_X1 port map( A1 => N4391, A2 => n16368, ZN => n16426);
   U15182 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n5368, ZN => n5740);
   U15183 : OAI221_X1 port map( B1 => n5747, B2 => n16361, C1 => n10385, C2 => 
                           n16362, A => n16427, ZN => n10450);
   U15184 : NAND2_X1 port map( A1 => N4496, A2 => n16364, ZN => n16427);
   U15185 : OAI221_X1 port map( B1 => n5747, B2 => n16365, C1 => n10353, C2 => 
                           n16366, A => n16428, ZN => n10449);
   U15186 : NAND2_X1 port map( A1 => N4390, A2 => n16368, ZN => n16428);
   U15187 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n5368, ZN => n5747);
   U15188 : OAI221_X1 port map( B1 => n5754, B2 => n16361, C1 => n10386, C2 => 
                           n16362, A => n16429, ZN => n10447);
   U15189 : NAND2_X1 port map( A1 => N4495, A2 => n16364, ZN => n16429);
   U15190 : OAI21_X1 port map( B1 => n16431, B2 => n16432, A => n16362, ZN => 
                           n16430);
   U15191 : INV_X1 port map( A => n16431, ZN => n16433);
   U15192 : NAND4_X1 port map( A1 => n16434, A2 => n16435, A3 => n16436, A4 => 
                           n16437, ZN => n16431);
   U15193 : NOR3_X1 port map( A1 => n16438, A2 => n16439, A3 => n16440, ZN => 
                           n16437);
   U15194 : XNOR2_X1 port map( A => r3013_A_4_port, B => n8743, ZN => n16440);
   U15195 : XNOR2_X1 port map( A => n581, B => n10076, ZN => n16439);
   U15196 : AND2_X1 port map( A1 => n16441, A2 => N3582, ZN => r3013_A_2_port);
   U15197 : XNOR2_X1 port map( A => r3013_A_3_port, B => n8742, ZN => n16438);
   U15198 : XNOR2_X1 port map( A => n10225, B => n646, ZN => n16436);
   U15199 : MUX2_X1 port map( A => RD2_ADD(0), B => N3580, S => n16441, Z => 
                           r3013_A_0_port);
   U15200 : XOR2_X1 port map( A => n6376, B => ADD_RD2_5_port, Z => n16435);
   U15201 : XNOR2_X1 port map( A => n11857, B => n594, ZN => n16434);
   U15202 : MUX2_X1 port map( A => RD2_ADD(1), B => N3581, S => n16441, Z => 
                           r3013_A_1_port);
   U15203 : OAI221_X1 port map( B1 => n5754, B2 => n16365, C1 => n10354, C2 => 
                           n16366, A => n16442, ZN => n10446);
   U15204 : NAND2_X1 port map( A1 => N4389, A2 => n16368, ZN => n16442);
   U15205 : OAI21_X1 port map( B1 => n16432, B2 => n16444, A => n16366, ZN => 
                           n16443);
   U15206 : NAND2_X1 port map( A1 => WR, A2 => n5368, ZN => n16432);
   U15207 : INV_X1 port map( A => n16444, ZN => n16445);
   U15208 : NAND4_X1 port map( A1 => n16446, A2 => n16447, A3 => n16448, A4 => 
                           n16449, ZN => n16444);
   U15209 : NOR3_X1 port map( A1 => n16450, A2 => n16451, A3 => n16452, ZN => 
                           n16449);
   U15210 : XNOR2_X1 port map( A => r3007_A_4_port, B => n8743, ZN => n16452);
   U15211 : NAND2_X1 port map( A1 => n16453, A2 => N3597, ZN => n8743);
   U15212 : XNOR2_X1 port map( A => ADD_RD1_5_port, B => n6376, ZN => n16451);
   U15213 : NAND2_X1 port map( A1 => N3598, A2 => n16453, ZN => n6376);
   U15214 : XNOR2_X1 port map( A => r3007_A_3_port, B => n8742, ZN => n16450);
   U15215 : NAND2_X1 port map( A1 => n16453, A2 => N3596, ZN => n8742);
   U15216 : XNOR2_X1 port map( A => n11857, B => n680, ZN => n16448);
   U15217 : MUX2_X1 port map( A => RD1_ADD(1), B => N3568, S => n16454, Z => 
                           r3007_A_1_port);
   U15218 : MUX2_X1 port map( A => WR_ADD(1), B => N3594, S => n16453, Z => 
                           n11857);
   U15219 : XNOR2_X1 port map( A => n10225, B => n732, ZN => n16447);
   U15220 : MUX2_X1 port map( A => RD1_ADD(0), B => N3567, S => n16454, Z => 
                           r3007_A_0_port);
   U15221 : MUX2_X1 port map( A => WR_ADD(0), B => N3593, S => n16453, Z => 
                           n10225);
   U15222 : XOR2_X1 port map( A => n10076, B => n668, Z => n16446);
   U15223 : AND2_X1 port map( A1 => n16454, A2 => N3569, ZN => r3007_A_2_port);
   U15224 : NAND2_X1 port map( A1 => n16453, A2 => N3595, ZN => n10076);
   U15225 : OR3_X1 port map( A1 => WR_ADD(4), A2 => WR_ADD(3), A3 => WR_ADD(2),
                           ZN => n16453);
   U15226 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n5368, ZN => n5754);
   U15227 : INV_X1 port map( A => WR_ADD(2), ZN => N3590);
   U15228 : INV_X1 port map( A => RD2_ADD(2), ZN => N3577);
   U15229 : INV_X1 port map( A => RD1_ADD(2), ZN => N3564);
   U15230 : OR3_X1 port map( A1 => RD2_ADD(4), A2 => RD2_ADD(3), A3 => 
                           RD2_ADD(2), ZN => n16441);
   U15231 : OR3_X1 port map( A1 => RD1_ADD(4), A2 => RD1_ADD(3), A3 => 
                           RD1_ADD(2), ZN => n16454);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N5_0 is

   port( a, b : in std_logic_vector (4 downto 0);  sel : in std_logic;  y : out
         std_logic_vector (4 downto 0));

end MUX21_N5_0;

architecture SYN_beh of MUX21_N5_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));
   U2 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U3 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U4 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U5 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity OR_GATE is

   port( x, y : in std_logic;  z : out std_logic);

end OR_GATE;

architecture SYN_DF of OR_GATE is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => x, A2 => y, ZN => z);

end SYN_DF;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity adder_generic_nbit32 is

   port( a, b : in std_logic_vector (31 downto 0);  y : out std_logic_vector 
         (31 downto 0));

end adder_generic_nbit32;

architecture SYN_Behavioral of adder_generic_nbit32 is

   component adder_generic_nbit32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1511 : std_logic;

begin
   
   n1 <= '0';
   add_21 : adder_generic_nbit32_DW01_add_0 port map( A(31) => a(31), A(30) => 
                           a(30), A(29) => a(29), A(28) => a(28), A(27) => 
                           a(27), A(26) => a(26), A(25) => a(25), A(24) => 
                           a(24), A(23) => a(23), A(22) => a(22), A(21) => 
                           a(21), A(20) => a(20), A(19) => a(19), A(18) => 
                           a(18), A(17) => a(17), A(16) => a(16), A(15) => 
                           a(15), A(14) => a(14), A(13) => a(13), A(12) => 
                           a(12), A(11) => a(11), A(10) => a(10), A(9) => a(9),
                           A(8) => a(8), A(7) => a(7), A(6) => a(6), A(5) => 
                           a(5), A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1)
                           => a(1), A(0) => a(0), B(31) => b(31), B(30) => 
                           b(30), B(29) => b(29), B(28) => b(28), B(27) => 
                           b(27), B(26) => b(26), B(25) => b(25), B(24) => 
                           b(24), B(23) => b(23), B(22) => b(22), B(21) => 
                           b(21), B(20) => b(20), B(19) => b(19), B(18) => 
                           b(18), B(17) => b(17), B(16) => b(16), B(15) => 
                           b(15), B(14) => b(14), B(13) => b(13), B(12) => 
                           b(12), B(11) => b(11), B(10) => b(10), B(9) => b(9),
                           B(8) => b(8), B(7) => b(7), B(6) => b(6), B(5) => 
                           b(5), B(4) => b(4), B(3) => b(3), B(2) => b(2), B(1)
                           => b(1), B(0) => b(0), CI => n1, SUM(31) => y(31), 
                           SUM(30) => y(30), SUM(29) => y(29), SUM(28) => y(28)
                           , SUM(27) => y(27), SUM(26) => y(26), SUM(25) => 
                           y(25), SUM(24) => y(24), SUM(23) => y(23), SUM(22) 
                           => y(22), SUM(21) => y(21), SUM(20) => y(20), 
                           SUM(19) => y(19), SUM(18) => y(18), SUM(17) => y(17)
                           , SUM(16) => y(16), SUM(15) => y(15), SUM(14) => 
                           y(14), SUM(13) => y(13), SUM(12) => y(12), SUM(11) 
                           => y(11), SUM(10) => y(10), SUM(9) => y(9), SUM(8) 
                           => y(8), SUM(7) => y(7), SUM(6) => y(6), SUM(5) => 
                           y(5), SUM(4) => y(4), SUM(3) => y(3), SUM(2) => y(2)
                           , SUM(1) => y(1), SUM(0) => y(0), CO => n_1511);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity sign_ext is

   port( a : in std_logic_vector (31 downto 0);  s : in std_logic;  y : out 
         std_logic_vector (31 downto 0));

end sign_ext;

architecture SYN_Behavioral of sign_ext is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal y_31_port, N23, N24, N25, N26, N27, N28, N29, N30, N31, N33, n3, n1, 
      n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   y <= ( y_31_port, N33, N33, N33, N33, N33, N33, N31, N30, N29, N28, N27, N26
      , N25, N24, N23, a(15), a(14), a(13), a(12), a(11), a(10), a(9), a(8), 
      a(7), a(6), a(5), a(4), a(3), a(2), a(1), a(0) );
   
   y_reg_31_inst : DLH_X1 port map( G => n3, D => N33, Q => y_31_port);
   n3 <= '1';
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => N33);
   U4 : NAND2_X1 port map( A1 => s, A2 => a(25), ZN => n2);
   U5 : NAND2_X1 port map( A1 => n1, A2 => n4, ZN => N31);
   U6 : NAND2_X1 port map( A1 => a(24), A2 => s, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n1, A2 => n5, ZN => N30);
   U8 : NAND2_X1 port map( A1 => a(23), A2 => s, ZN => n5);
   U9 : NAND2_X1 port map( A1 => n1, A2 => n6, ZN => N29);
   U10 : NAND2_X1 port map( A1 => a(22), A2 => s, ZN => n6);
   U11 : NAND2_X1 port map( A1 => n1, A2 => n7, ZN => N28);
   U12 : NAND2_X1 port map( A1 => a(21), A2 => s, ZN => n7);
   U13 : NAND2_X1 port map( A1 => n1, A2 => n8, ZN => N27);
   U14 : NAND2_X1 port map( A1 => a(20), A2 => s, ZN => n8);
   U15 : NAND2_X1 port map( A1 => n1, A2 => n9, ZN => N26);
   U16 : NAND2_X1 port map( A1 => a(19), A2 => s, ZN => n9);
   U17 : NAND2_X1 port map( A1 => n1, A2 => n10, ZN => N25);
   U18 : NAND2_X1 port map( A1 => a(18), A2 => s, ZN => n10);
   U19 : NAND2_X1 port map( A1 => n1, A2 => n11, ZN => N24);
   U20 : NAND2_X1 port map( A1 => a(17), A2 => s, ZN => n11);
   U21 : NAND2_X1 port map( A1 => n1, A2 => n12, ZN => N23);
   U22 : NAND2_X1 port map( A1 => a(16), A2 => s, ZN => n12);
   U23 : NAND2_X1 port map( A1 => a(15), A2 => n13, ZN => n1);
   U24 : INV_X1 port map( A => s, ZN => n13);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity adder_genericu_nbit32 is

   port( a, b : in std_logic_vector (31 downto 0);  y : out std_logic_vector 
         (31 downto 0));

end adder_genericu_nbit32;

architecture SYN_Behavioral of adder_genericu_nbit32 is

   component adder_genericu_nbit32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1512 : std_logic;

begin
   
   n1 <= '0';
   add_13 : adder_genericu_nbit32_DW01_add_0 port map( A(31) => a(31), A(30) =>
                           a(30), A(29) => a(29), A(28) => a(28), A(27) => 
                           a(27), A(26) => a(26), A(25) => a(25), A(24) => 
                           a(24), A(23) => a(23), A(22) => a(22), A(21) => 
                           a(21), A(20) => a(20), A(19) => a(19), A(18) => 
                           a(18), A(17) => a(17), A(16) => a(16), A(15) => 
                           a(15), A(14) => a(14), A(13) => a(13), A(12) => 
                           a(12), A(11) => a(11), A(10) => a(10), A(9) => a(9),
                           A(8) => a(8), A(7) => a(7), A(6) => a(6), A(5) => 
                           a(5), A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1)
                           => a(1), A(0) => a(0), B(31) => b(31), B(30) => 
                           b(30), B(29) => b(29), B(28) => b(28), B(27) => 
                           b(27), B(26) => b(26), B(25) => b(25), B(24) => 
                           b(24), B(23) => b(23), B(22) => b(22), B(21) => 
                           b(21), B(20) => b(20), B(19) => b(19), B(18) => 
                           b(18), B(17) => b(17), B(16) => b(16), B(15) => 
                           b(15), B(14) => b(14), B(13) => b(13), B(12) => 
                           b(12), B(11) => b(11), B(10) => b(10), B(9) => b(9),
                           B(8) => b(8), B(7) => b(7), B(6) => b(6), B(5) => 
                           b(5), B(4) => b(4), B(3) => b(3), B(2) => b(2), B(1)
                           => b(1), B(0) => b(0), CI => n1, SUM(31) => y(31), 
                           SUM(30) => y(30), SUM(29) => y(29), SUM(28) => y(28)
                           , SUM(27) => y(27), SUM(26) => y(26), SUM(25) => 
                           y(25), SUM(24) => y(24), SUM(23) => y(23), SUM(22) 
                           => y(22), SUM(21) => y(21), SUM(20) => y(20), 
                           SUM(19) => y(19), SUM(18) => y(18), SUM(17) => y(17)
                           , SUM(16) => y(16), SUM(15) => y(15), SUM(14) => 
                           y(14), SUM(13) => y(13), SUM(12) => y(12), SUM(11) 
                           => y(11), SUM(10) => y(10), SUM(9) => y(9), SUM(8) 
                           => y(8), SUM(7) => y(7), SUM(6) => y(6), SUM(5) => 
                           y(5), SUM(4) => y(4), SUM(3) => y(3), SUM(2) => y(2)
                           , SUM(1) => y(1), SUM(0) => y(0), CO => n_1512);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity register_generic_nbit32 is

   port( d : in std_logic_vector (31 downto 0);  q : out std_logic_vector (31 
         downto 0);  clk, reset, en : in std_logic);

end register_generic_nbit32;

architecture SYN_Behavioral of register_generic_nbit32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal q_31_port, q_30_port, q_29_port, q_28_port, q_27_port, q_26_port, 
      q_25_port, q_24_port, q_23_port, q_22_port, q_21_port, q_20_port, 
      q_19_port, q_18_port, q_17_port, q_16_port, q_15_port, q_14_port, 
      q_13_port, q_12_port, q_11_port, q_10_port, q_9_port, q_8_port, q_7_port,
      q_6_port, q_5_port, q_4_port, q_3_port, q_2_port, q_1_port, q_0_port, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n97, n1, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544 : std_logic;

begin
   q <= ( q_31_port, q_30_port, q_29_port, q_28_port, q_27_port, q_26_port, 
      q_25_port, q_24_port, q_23_port, q_22_port, q_21_port, q_20_port, 
      q_19_port, q_18_port, q_17_port, q_16_port, q_15_port, q_14_port, 
      q_13_port, q_12_port, q_11_port, q_10_port, q_9_port, q_8_port, q_7_port,
      q_6_port, q_5_port, q_4_port, q_3_port, q_2_port, q_1_port, q_0_port );
   
   q_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n1, Q => 
                           q_31_port, QN => n_1513);
   q_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n1, Q => 
                           q_30_port, QN => n_1514);
   q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n1, Q => 
                           q_29_port, QN => n_1515);
   q_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n1, Q => 
                           q_28_port, QN => n_1516);
   q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n1, Q => 
                           q_27_port, QN => n_1517);
   q_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n1, Q => 
                           q_26_port, QN => n_1518);
   q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n1, Q => 
                           q_25_port, QN => n_1519);
   q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n1, Q => 
                           q_24_port, QN => n_1520);
   q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n1, Q => 
                           q_23_port, QN => n_1521);
   q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n1, Q => 
                           q_22_port, QN => n_1522);
   q_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n1, Q => 
                           q_21_port, QN => n_1523);
   q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n1, Q => 
                           q_20_port, QN => n_1524);
   q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n1, Q => 
                           q_19_port, QN => n_1525);
   q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n1, Q => 
                           q_18_port, QN => n_1526);
   q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n1, Q => 
                           q_17_port, QN => n_1527);
   q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n1, Q => 
                           q_16_port, QN => n_1528);
   q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n1, Q => 
                           q_15_port, QN => n_1529);
   q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n1, Q => 
                           q_14_port, QN => n_1530);
   q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n1, Q => 
                           q_13_port, QN => n_1531);
   q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n1, Q => 
                           q_12_port, QN => n_1532);
   q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n1, Q => 
                           q_11_port, QN => n_1533);
   q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n1, Q => 
                           q_10_port, QN => n_1534);
   q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n1, Q => 
                           q_9_port, QN => n_1535);
   q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n1, Q => 
                           q_8_port, QN => n_1536);
   q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n1, Q => 
                           q_7_port, QN => n_1537);
   q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n1, Q => 
                           q_6_port, QN => n_1538);
   q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n1, Q => 
                           q_5_port, QN => n_1539);
   q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n1, Q => 
                           q_4_port, QN => n_1540);
   q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n1, Q => 
                           q_3_port, QN => n_1541);
   q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n1, Q => 
                           q_2_port, QN => n_1542);
   q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n1, Q => 
                           q_1_port, QN => n_1543);
   q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n1, Q => 
                           q_0_port, QN => n_1544);
   U2 : INV_X2 port map( A => reset, ZN => n1);
   U3 : MUX2_X1 port map( A => q_31_port, B => d(31), S => en, Z => n97);
   U4 : MUX2_X1 port map( A => q_30_port, B => d(30), S => en, Z => n95);
   U5 : MUX2_X1 port map( A => q_29_port, B => d(29), S => en, Z => n94);
   U6 : MUX2_X1 port map( A => q_28_port, B => d(28), S => en, Z => n93);
   U7 : MUX2_X1 port map( A => q_27_port, B => d(27), S => en, Z => n92);
   U8 : MUX2_X1 port map( A => q_26_port, B => d(26), S => en, Z => n91);
   U9 : MUX2_X1 port map( A => q_25_port, B => d(25), S => en, Z => n90);
   U10 : MUX2_X1 port map( A => q_24_port, B => d(24), S => en, Z => n89);
   U11 : MUX2_X1 port map( A => q_23_port, B => d(23), S => en, Z => n88);
   U12 : MUX2_X1 port map( A => q_22_port, B => d(22), S => en, Z => n87);
   U13 : MUX2_X1 port map( A => q_21_port, B => d(21), S => en, Z => n86);
   U14 : MUX2_X1 port map( A => q_20_port, B => d(20), S => en, Z => n85);
   U15 : MUX2_X1 port map( A => q_19_port, B => d(19), S => en, Z => n84);
   U16 : MUX2_X1 port map( A => q_18_port, B => d(18), S => en, Z => n83);
   U17 : MUX2_X1 port map( A => q_17_port, B => d(17), S => en, Z => n82);
   U18 : MUX2_X1 port map( A => q_16_port, B => d(16), S => en, Z => n81);
   U19 : MUX2_X1 port map( A => q_15_port, B => d(15), S => en, Z => n80);
   U20 : MUX2_X1 port map( A => q_14_port, B => d(14), S => en, Z => n79);
   U21 : MUX2_X1 port map( A => q_13_port, B => d(13), S => en, Z => n78);
   U22 : MUX2_X1 port map( A => q_12_port, B => d(12), S => en, Z => n77);
   U23 : MUX2_X1 port map( A => q_11_port, B => d(11), S => en, Z => n76);
   U24 : MUX2_X1 port map( A => q_10_port, B => d(10), S => en, Z => n75);
   U25 : MUX2_X1 port map( A => q_9_port, B => d(9), S => en, Z => n74);
   U26 : MUX2_X1 port map( A => q_8_port, B => d(8), S => en, Z => n73);
   U27 : MUX2_X1 port map( A => q_7_port, B => d(7), S => en, Z => n72);
   U28 : MUX2_X1 port map( A => q_6_port, B => d(6), S => en, Z => n71);
   U29 : MUX2_X1 port map( A => q_5_port, B => d(5), S => en, Z => n70);
   U30 : MUX2_X1 port map( A => q_4_port, B => d(4), S => en, Z => n69);
   U31 : MUX2_X1 port map( A => q_3_port, B => d(3), S => en, Z => n68);
   U32 : MUX2_X1 port map( A => q_2_port, B => d(2), S => en, Z => n67);
   U33 : MUX2_X1 port map( A => q_1_port, B => d(1), S => en, Z => n66);
   U34 : MUX2_X1 port map( A => q_0_port, B => d(0), S => en, Z => n65);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity MUX21_N32_0 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end MUX21_N32_0;

architecture SYN_beh of MUX21_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => a(31), B => b(31), S => sel, Z => y(31));
   U2 : MUX2_X1 port map( A => a(30), B => b(30), S => sel, Z => y(30));
   U3 : MUX2_X1 port map( A => a(29), B => b(29), S => sel, Z => y(29));
   U4 : MUX2_X1 port map( A => a(28), B => b(28), S => sel, Z => y(28));
   U5 : MUX2_X1 port map( A => a(27), B => b(27), S => sel, Z => y(27));
   U6 : MUX2_X1 port map( A => a(26), B => b(26), S => sel, Z => y(26));
   U7 : MUX2_X1 port map( A => a(25), B => b(25), S => sel, Z => y(25));
   U8 : MUX2_X1 port map( A => a(24), B => b(24), S => sel, Z => y(24));
   U9 : MUX2_X1 port map( A => a(23), B => b(23), S => sel, Z => y(23));
   U10 : MUX2_X1 port map( A => a(22), B => b(22), S => sel, Z => y(22));
   U11 : MUX2_X1 port map( A => a(21), B => b(21), S => sel, Z => y(21));
   U12 : MUX2_X1 port map( A => a(20), B => b(20), S => sel, Z => y(20));
   U13 : MUX2_X1 port map( A => a(19), B => b(19), S => sel, Z => y(19));
   U14 : MUX2_X1 port map( A => a(18), B => b(18), S => sel, Z => y(18));
   U15 : MUX2_X1 port map( A => a(17), B => b(17), S => sel, Z => y(17));
   U16 : MUX2_X1 port map( A => a(16), B => b(16), S => sel, Z => y(16));
   U17 : MUX2_X1 port map( A => a(15), B => b(15), S => sel, Z => y(15));
   U18 : MUX2_X1 port map( A => a(14), B => b(14), S => sel, Z => y(14));
   U19 : MUX2_X1 port map( A => a(13), B => b(13), S => sel, Z => y(13));
   U20 : MUX2_X1 port map( A => a(12), B => b(12), S => sel, Z => y(12));
   U21 : MUX2_X1 port map( A => a(11), B => b(11), S => sel, Z => y(11));
   U22 : MUX2_X1 port map( A => a(10), B => b(10), S => sel, Z => y(10));
   U23 : MUX2_X1 port map( A => a(9), B => b(9), S => sel, Z => y(9));
   U24 : MUX2_X1 port map( A => a(8), B => b(8), S => sel, Z => y(8));
   U25 : MUX2_X1 port map( A => a(7), B => b(7), S => sel, Z => y(7));
   U26 : MUX2_X1 port map( A => a(6), B => b(6), S => sel, Z => y(6));
   U27 : MUX2_X1 port map( A => a(5), B => b(5), S => sel, Z => y(5));
   U28 : MUX2_X1 port map( A => a(4), B => b(4), S => sel, Z => y(4));
   U29 : MUX2_X1 port map( A => a(3), B => b(3), S => sel, Z => y(3));
   U30 : MUX2_X1 port map( A => a(2), B => b(2), S => sel, Z => y(2));
   U31 : MUX2_X1 port map( A => a(1), B => b(1), S => sel, Z => y(1));
   U32 : MUX2_X1 port map( A => a(0), B => b(0), S => sel, Z => y(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity writeback_unit_N32 is

   port( ReadDataW, ALUOutW : in std_logic_vector (31 downto 0);  WriteRegW : 
         in std_logic_vector (4 downto 0);  MemToRegW : in std_logic;  
         WriteRegW_out : out std_logic_vector (4 downto 0);  ResultW : out 
         std_logic_vector (31 downto 0));

end writeback_unit_N32;

architecture SYN_Structural of writeback_unit_N32 is

   component MUX21_N32_2
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;

begin
   WriteRegW_out <= ( WriteRegW(4), WriteRegW(3), WriteRegW(2), WriteRegW(1), 
      WriteRegW(0) );
   
   MUX21_1 : MUX21_N32_2 port map( a(31) => ALUOutW(31), a(30) => ALUOutW(30), 
                           a(29) => ALUOutW(29), a(28) => ALUOutW(28), a(27) =>
                           ALUOutW(27), a(26) => ALUOutW(26), a(25) => 
                           ALUOutW(25), a(24) => ALUOutW(24), a(23) => 
                           ALUOutW(23), a(22) => ALUOutW(22), a(21) => 
                           ALUOutW(21), a(20) => ALUOutW(20), a(19) => 
                           ALUOutW(19), a(18) => ALUOutW(18), a(17) => 
                           ALUOutW(17), a(16) => ALUOutW(16), a(15) => 
                           ALUOutW(15), a(14) => ALUOutW(14), a(13) => 
                           ALUOutW(13), a(12) => ALUOutW(12), a(11) => 
                           ALUOutW(11), a(10) => ALUOutW(10), a(9) => 
                           ALUOutW(9), a(8) => ALUOutW(8), a(7) => ALUOutW(7), 
                           a(6) => ALUOutW(6), a(5) => ALUOutW(5), a(4) => 
                           ALUOutW(4), a(3) => ALUOutW(3), a(2) => ALUOutW(2), 
                           a(1) => ALUOutW(1), a(0) => ALUOutW(0), b(31) => 
                           ReadDataW(31), b(30) => ReadDataW(30), b(29) => 
                           ReadDataW(29), b(28) => ReadDataW(28), b(27) => 
                           ReadDataW(27), b(26) => ReadDataW(26), b(25) => 
                           ReadDataW(25), b(24) => ReadDataW(24), b(23) => 
                           ReadDataW(23), b(22) => ReadDataW(22), b(21) => 
                           ReadDataW(21), b(20) => ReadDataW(20), b(19) => 
                           ReadDataW(19), b(18) => ReadDataW(18), b(17) => 
                           ReadDataW(17), b(16) => ReadDataW(16), b(15) => 
                           ReadDataW(15), b(14) => ReadDataW(14), b(13) => 
                           ReadDataW(13), b(12) => ReadDataW(12), b(11) => 
                           ReadDataW(11), b(10) => ReadDataW(10), b(9) => 
                           ReadDataW(9), b(8) => ReadDataW(8), b(7) => 
                           ReadDataW(7), b(6) => ReadDataW(6), b(5) => 
                           ReadDataW(5), b(4) => ReadDataW(4), b(3) => 
                           ReadDataW(3), b(2) => ReadDataW(2), b(1) => 
                           ReadDataW(1), b(0) => ReadDataW(0), sel => MemToRegW
                           , y(31) => ResultW(31), y(30) => ResultW(30), y(29) 
                           => ResultW(29), y(28) => ResultW(28), y(27) => 
                           ResultW(27), y(26) => ResultW(26), y(25) => 
                           ResultW(25), y(24) => ResultW(24), y(23) => 
                           ResultW(23), y(22) => ResultW(22), y(21) => 
                           ResultW(21), y(20) => ResultW(20), y(19) => 
                           ResultW(19), y(18) => ResultW(18), y(17) => 
                           ResultW(17), y(16) => ResultW(16), y(15) => 
                           ResultW(15), y(14) => ResultW(14), y(13) => 
                           ResultW(13), y(12) => ResultW(12), y(11) => 
                           ResultW(11), y(10) => ResultW(10), y(9) => 
                           ResultW(9), y(8) => ResultW(8), y(7) => ResultW(7), 
                           y(6) => ResultW(6), y(5) => ResultW(5), y(4) => 
                           ResultW(4), y(3) => ResultW(3), y(2) => ResultW(2), 
                           y(1) => ResultW(1), y(0) => ResultW(0));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity memory_unit_nbit32_nwords64 is

   port( ALUOutMIn, WriteDataM : in std_logic_vector (31 downto 0);  ReadDataM,
         ALUOutMOut, address_to_dram, data_to_dram : out std_logic_vector (31 
         downto 0);  dram_to_dlx : in std_logic_vector (31 downto 0);  
         WriteRegMIn : in std_logic_vector (4 downto 0);  WriteRegMOut : out 
         std_logic_vector (4 downto 0);  clk, rst, MemWriteM : in std_logic;  
         MemWriteM_out : out std_logic);

end memory_unit_nbit32_nwords64;

architecture SYN_Structural of memory_unit_nbit32_nwords64 is

begin
   ReadDataM <= ( dram_to_dlx(31), dram_to_dlx(30), dram_to_dlx(29), 
      dram_to_dlx(28), dram_to_dlx(27), dram_to_dlx(26), dram_to_dlx(25), 
      dram_to_dlx(24), dram_to_dlx(23), dram_to_dlx(22), dram_to_dlx(21), 
      dram_to_dlx(20), dram_to_dlx(19), dram_to_dlx(18), dram_to_dlx(17), 
      dram_to_dlx(16), dram_to_dlx(15), dram_to_dlx(14), dram_to_dlx(13), 
      dram_to_dlx(12), dram_to_dlx(11), dram_to_dlx(10), dram_to_dlx(9), 
      dram_to_dlx(8), dram_to_dlx(7), dram_to_dlx(6), dram_to_dlx(5), 
      dram_to_dlx(4), dram_to_dlx(3), dram_to_dlx(2), dram_to_dlx(1), 
      dram_to_dlx(0) );
   ALUOutMOut <= ( ALUOutMIn(31), ALUOutMIn(30), ALUOutMIn(29), ALUOutMIn(28), 
      ALUOutMIn(27), ALUOutMIn(26), ALUOutMIn(25), ALUOutMIn(24), ALUOutMIn(23)
      , ALUOutMIn(22), ALUOutMIn(21), ALUOutMIn(20), ALUOutMIn(19), 
      ALUOutMIn(18), ALUOutMIn(17), ALUOutMIn(16), ALUOutMIn(15), ALUOutMIn(14)
      , ALUOutMIn(13), ALUOutMIn(12), ALUOutMIn(11), ALUOutMIn(10), 
      ALUOutMIn(9), ALUOutMIn(8), ALUOutMIn(7), ALUOutMIn(6), ALUOutMIn(5), 
      ALUOutMIn(4), ALUOutMIn(3), ALUOutMIn(2), ALUOutMIn(1), ALUOutMIn(0) );
   address_to_dram <= ( ALUOutMIn(31), ALUOutMIn(30), ALUOutMIn(29), 
      ALUOutMIn(28), ALUOutMIn(27), ALUOutMIn(26), ALUOutMIn(25), ALUOutMIn(24)
      , ALUOutMIn(23), ALUOutMIn(22), ALUOutMIn(21), ALUOutMIn(20), 
      ALUOutMIn(19), ALUOutMIn(18), ALUOutMIn(17), ALUOutMIn(16), ALUOutMIn(15)
      , ALUOutMIn(14), ALUOutMIn(13), ALUOutMIn(12), ALUOutMIn(11), 
      ALUOutMIn(10), ALUOutMIn(9), ALUOutMIn(8), ALUOutMIn(7), ALUOutMIn(6), 
      ALUOutMIn(5), ALUOutMIn(4), ALUOutMIn(3), ALUOutMIn(2), ALUOutMIn(1), 
      ALUOutMIn(0) );
   data_to_dram <= ( WriteDataM(31), WriteDataM(30), WriteDataM(29), 
      WriteDataM(28), WriteDataM(27), WriteDataM(26), WriteDataM(25), 
      WriteDataM(24), WriteDataM(23), WriteDataM(22), WriteDataM(21), 
      WriteDataM(20), WriteDataM(19), WriteDataM(18), WriteDataM(17), 
      WriteDataM(16), WriteDataM(15), WriteDataM(14), WriteDataM(13), 
      WriteDataM(12), WriteDataM(11), WriteDataM(10), WriteDataM(9), 
      WriteDataM(8), WriteDataM(7), WriteDataM(6), WriteDataM(5), WriteDataM(4)
      , WriteDataM(3), WriteDataM(2), WriteDataM(1), WriteDataM(0) );
   WriteRegMOut <= ( WriteRegMIn(4), WriteRegMIn(3), WriteRegMIn(2), 
      WriteRegMIn(1), WriteRegMIn(0) );
   MemWriteM_out <= MemWriteM;

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity execute_stage_wrapper_NBIT32_N32 is

   port( en_alu : in std_logic;  RD1E, RD2E : in std_logic_vector (31 downto 0)
         ;  RsE, RdE, RtE : in std_logic_vector (4 downto 0);  SignImmE, 
         ALUOutME, ResultWE : in std_logic_vector (31 downto 0);  ALUoutE : out
         std_logic_vector (31 downto 0);  WriteRegE : out std_logic_vector (4 
         downto 0);  WriteDataE : out std_logic_vector (31 downto 0);  
         ForwardAE, ForwardBE : in std_logic_vector (1 downto 0);  RsE_o, RtE_o
         : out std_logic_vector (4 downto 0);  RegDstE, ALUSrcE : in std_logic;
         ALUcontrolE : in std_logic_vector (5 downto 0));

end execute_stage_wrapper_NBIT32_N32;

architecture SYN_Behavioral of execute_stage_wrapper_NBIT32_N32 is

   component ALU_NBIT32
      port( en_alu : in std_logic;  op1, op2 : in std_logic_vector (31 downto 
            0);  sel : in std_logic_vector (5 downto 0);  result : out 
            std_logic_vector (31 downto 0);  CarryOut, overflow : out std_logic
            );
   end component;
   
   component MUX21_N5_1
      port( a, b : in std_logic_vector (4 downto 0);  sel : in std_logic;  y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX21_N32_3
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux31_N32_1
      port( a, b, c : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  y : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux31_N32_0
      port( a, b, c : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  y : out std_logic_vector (31 downto
            0));
   end component;
   
   signal WriteDataE_31_port, WriteDataE_30_port, WriteDataE_29_port, 
      WriteDataE_28_port, WriteDataE_27_port, WriteDataE_26_port, 
      WriteDataE_25_port, WriteDataE_24_port, WriteDataE_23_port, 
      WriteDataE_22_port, WriteDataE_21_port, WriteDataE_20_port, 
      WriteDataE_19_port, WriteDataE_18_port, WriteDataE_17_port, 
      WriteDataE_16_port, WriteDataE_15_port, WriteDataE_14_port, 
      WriteDataE_13_port, WriteDataE_12_port, WriteDataE_11_port, 
      WriteDataE_10_port, WriteDataE_9_port, WriteDataE_8_port, 
      WriteDataE_7_port, WriteDataE_6_port, WriteDataE_5_port, 
      WriteDataE_4_port, WriteDataE_3_port, WriteDataE_2_port, 
      WriteDataE_1_port, WriteDataE_0_port, SrcAE_31_port, SrcAE_30_port, 
      SrcAE_29_port, SrcAE_28_port, SrcAE_27_port, SrcAE_26_port, SrcAE_25_port
      , SrcAE_24_port, SrcAE_23_port, SrcAE_22_port, SrcAE_21_port, 
      SrcAE_20_port, SrcAE_19_port, SrcAE_18_port, SrcAE_17_port, SrcAE_16_port
      , SrcAE_15_port, SrcAE_14_port, SrcAE_13_port, SrcAE_12_port, 
      SrcAE_11_port, SrcAE_10_port, SrcAE_9_port, SrcAE_8_port, SrcAE_7_port, 
      SrcAE_6_port, SrcAE_5_port, SrcAE_4_port, SrcAE_3_port, SrcAE_2_port, 
      SrcAE_1_port, SrcAE_0_port, SrcBE_31_port, SrcBE_30_port, SrcBE_29_port, 
      SrcBE_28_port, SrcBE_27_port, SrcBE_26_port, SrcBE_25_port, SrcBE_24_port
      , SrcBE_23_port, SrcBE_22_port, SrcBE_21_port, SrcBE_20_port, 
      SrcBE_19_port, SrcBE_18_port, SrcBE_17_port, SrcBE_16_port, SrcBE_15_port
      , SrcBE_14_port, SrcBE_13_port, SrcBE_12_port, SrcBE_11_port, 
      SrcBE_10_port, SrcBE_9_port, SrcBE_8_port, SrcBE_7_port, SrcBE_6_port, 
      SrcBE_5_port, SrcBE_4_port, SrcBE_3_port, SrcBE_2_port, SrcBE_1_port, 
      SrcBE_0_port, n_1545, n_1546 : std_logic;

begin
   WriteDataE <= ( WriteDataE_31_port, WriteDataE_30_port, WriteDataE_29_port, 
      WriteDataE_28_port, WriteDataE_27_port, WriteDataE_26_port, 
      WriteDataE_25_port, WriteDataE_24_port, WriteDataE_23_port, 
      WriteDataE_22_port, WriteDataE_21_port, WriteDataE_20_port, 
      WriteDataE_19_port, WriteDataE_18_port, WriteDataE_17_port, 
      WriteDataE_16_port, WriteDataE_15_port, WriteDataE_14_port, 
      WriteDataE_13_port, WriteDataE_12_port, WriteDataE_11_port, 
      WriteDataE_10_port, WriteDataE_9_port, WriteDataE_8_port, 
      WriteDataE_7_port, WriteDataE_6_port, WriteDataE_5_port, 
      WriteDataE_4_port, WriteDataE_3_port, WriteDataE_2_port, 
      WriteDataE_1_port, WriteDataE_0_port );
   RsE_o <= ( RsE(4), RsE(3), RsE(2), RsE(1), RsE(0) );
   RtE_o <= ( RtE(4), RtE(3), RtE(2), RtE(1), RtE(0) );
   
   mux31_1 : mux31_N32_0 port map( a(31) => RD1E(31), a(30) => RD1E(30), a(29) 
                           => RD1E(29), a(28) => RD1E(28), a(27) => RD1E(27), 
                           a(26) => RD1E(26), a(25) => RD1E(25), a(24) => 
                           RD1E(24), a(23) => RD1E(23), a(22) => RD1E(22), 
                           a(21) => RD1E(21), a(20) => RD1E(20), a(19) => 
                           RD1E(19), a(18) => RD1E(18), a(17) => RD1E(17), 
                           a(16) => RD1E(16), a(15) => RD1E(15), a(14) => 
                           RD1E(14), a(13) => RD1E(13), a(12) => RD1E(12), 
                           a(11) => RD1E(11), a(10) => RD1E(10), a(9) => 
                           RD1E(9), a(8) => RD1E(8), a(7) => RD1E(7), a(6) => 
                           RD1E(6), a(5) => RD1E(5), a(4) => RD1E(4), a(3) => 
                           RD1E(3), a(2) => RD1E(2), a(1) => RD1E(1), a(0) => 
                           RD1E(0), b(31) => ResultWE(31), b(30) => 
                           ResultWE(30), b(29) => ResultWE(29), b(28) => 
                           ResultWE(28), b(27) => ResultWE(27), b(26) => 
                           ResultWE(26), b(25) => ResultWE(25), b(24) => 
                           ResultWE(24), b(23) => ResultWE(23), b(22) => 
                           ResultWE(22), b(21) => ResultWE(21), b(20) => 
                           ResultWE(20), b(19) => ResultWE(19), b(18) => 
                           ResultWE(18), b(17) => ResultWE(17), b(16) => 
                           ResultWE(16), b(15) => ResultWE(15), b(14) => 
                           ResultWE(14), b(13) => ResultWE(13), b(12) => 
                           ResultWE(12), b(11) => ResultWE(11), b(10) => 
                           ResultWE(10), b(9) => ResultWE(9), b(8) => 
                           ResultWE(8), b(7) => ResultWE(7), b(6) => 
                           ResultWE(6), b(5) => ResultWE(5), b(4) => 
                           ResultWE(4), b(3) => ResultWE(3), b(2) => 
                           ResultWE(2), b(1) => ResultWE(1), b(0) => 
                           ResultWE(0), c(31) => ALUOutME(31), c(30) => 
                           ALUOutME(30), c(29) => ALUOutME(29), c(28) => 
                           ALUOutME(28), c(27) => ALUOutME(27), c(26) => 
                           ALUOutME(26), c(25) => ALUOutME(25), c(24) => 
                           ALUOutME(24), c(23) => ALUOutME(23), c(22) => 
                           ALUOutME(22), c(21) => ALUOutME(21), c(20) => 
                           ALUOutME(20), c(19) => ALUOutME(19), c(18) => 
                           ALUOutME(18), c(17) => ALUOutME(17), c(16) => 
                           ALUOutME(16), c(15) => ALUOutME(15), c(14) => 
                           ALUOutME(14), c(13) => ALUOutME(13), c(12) => 
                           ALUOutME(12), c(11) => ALUOutME(11), c(10) => 
                           ALUOutME(10), c(9) => ALUOutME(9), c(8) => 
                           ALUOutME(8), c(7) => ALUOutME(7), c(6) => 
                           ALUOutME(6), c(5) => ALUOutME(5), c(4) => 
                           ALUOutME(4), c(3) => ALUOutME(3), c(2) => 
                           ALUOutME(2), c(1) => ALUOutME(1), c(0) => 
                           ALUOutME(0), sel(1) => ForwardAE(1), sel(0) => 
                           ForwardAE(0), y(31) => SrcAE_31_port, y(30) => 
                           SrcAE_30_port, y(29) => SrcAE_29_port, y(28) => 
                           SrcAE_28_port, y(27) => SrcAE_27_port, y(26) => 
                           SrcAE_26_port, y(25) => SrcAE_25_port, y(24) => 
                           SrcAE_24_port, y(23) => SrcAE_23_port, y(22) => 
                           SrcAE_22_port, y(21) => SrcAE_21_port, y(20) => 
                           SrcAE_20_port, y(19) => SrcAE_19_port, y(18) => 
                           SrcAE_18_port, y(17) => SrcAE_17_port, y(16) => 
                           SrcAE_16_port, y(15) => SrcAE_15_port, y(14) => 
                           SrcAE_14_port, y(13) => SrcAE_13_port, y(12) => 
                           SrcAE_12_port, y(11) => SrcAE_11_port, y(10) => 
                           SrcAE_10_port, y(9) => SrcAE_9_port, y(8) => 
                           SrcAE_8_port, y(7) => SrcAE_7_port, y(6) => 
                           SrcAE_6_port, y(5) => SrcAE_5_port, y(4) => 
                           SrcAE_4_port, y(3) => SrcAE_3_port, y(2) => 
                           SrcAE_2_port, y(1) => SrcAE_1_port, y(0) => 
                           SrcAE_0_port);
   mex31_2 : mux31_N32_1 port map( a(31) => RD2E(31), a(30) => RD2E(30), a(29) 
                           => RD2E(29), a(28) => RD2E(28), a(27) => RD2E(27), 
                           a(26) => RD2E(26), a(25) => RD2E(25), a(24) => 
                           RD2E(24), a(23) => RD2E(23), a(22) => RD2E(22), 
                           a(21) => RD2E(21), a(20) => RD2E(20), a(19) => 
                           RD2E(19), a(18) => RD2E(18), a(17) => RD2E(17), 
                           a(16) => RD2E(16), a(15) => RD2E(15), a(14) => 
                           RD2E(14), a(13) => RD2E(13), a(12) => RD2E(12), 
                           a(11) => RD2E(11), a(10) => RD2E(10), a(9) => 
                           RD2E(9), a(8) => RD2E(8), a(7) => RD2E(7), a(6) => 
                           RD2E(6), a(5) => RD2E(5), a(4) => RD2E(4), a(3) => 
                           RD2E(3), a(2) => RD2E(2), a(1) => RD2E(1), a(0) => 
                           RD2E(0), b(31) => ResultWE(31), b(30) => 
                           ResultWE(30), b(29) => ResultWE(29), b(28) => 
                           ResultWE(28), b(27) => ResultWE(27), b(26) => 
                           ResultWE(26), b(25) => ResultWE(25), b(24) => 
                           ResultWE(24), b(23) => ResultWE(23), b(22) => 
                           ResultWE(22), b(21) => ResultWE(21), b(20) => 
                           ResultWE(20), b(19) => ResultWE(19), b(18) => 
                           ResultWE(18), b(17) => ResultWE(17), b(16) => 
                           ResultWE(16), b(15) => ResultWE(15), b(14) => 
                           ResultWE(14), b(13) => ResultWE(13), b(12) => 
                           ResultWE(12), b(11) => ResultWE(11), b(10) => 
                           ResultWE(10), b(9) => ResultWE(9), b(8) => 
                           ResultWE(8), b(7) => ResultWE(7), b(6) => 
                           ResultWE(6), b(5) => ResultWE(5), b(4) => 
                           ResultWE(4), b(3) => ResultWE(3), b(2) => 
                           ResultWE(2), b(1) => ResultWE(1), b(0) => 
                           ResultWE(0), c(31) => ALUOutME(31), c(30) => 
                           ALUOutME(30), c(29) => ALUOutME(29), c(28) => 
                           ALUOutME(28), c(27) => ALUOutME(27), c(26) => 
                           ALUOutME(26), c(25) => ALUOutME(25), c(24) => 
                           ALUOutME(24), c(23) => ALUOutME(23), c(22) => 
                           ALUOutME(22), c(21) => ALUOutME(21), c(20) => 
                           ALUOutME(20), c(19) => ALUOutME(19), c(18) => 
                           ALUOutME(18), c(17) => ALUOutME(17), c(16) => 
                           ALUOutME(16), c(15) => ALUOutME(15), c(14) => 
                           ALUOutME(14), c(13) => ALUOutME(13), c(12) => 
                           ALUOutME(12), c(11) => ALUOutME(11), c(10) => 
                           ALUOutME(10), c(9) => ALUOutME(9), c(8) => 
                           ALUOutME(8), c(7) => ALUOutME(7), c(6) => 
                           ALUOutME(6), c(5) => ALUOutME(5), c(4) => 
                           ALUOutME(4), c(3) => ALUOutME(3), c(2) => 
                           ALUOutME(2), c(1) => ALUOutME(1), c(0) => 
                           ALUOutME(0), sel(1) => ForwardBE(1), sel(0) => 
                           ForwardBE(0), y(31) => WriteDataE_31_port, y(30) => 
                           WriteDataE_30_port, y(29) => WriteDataE_29_port, 
                           y(28) => WriteDataE_28_port, y(27) => 
                           WriteDataE_27_port, y(26) => WriteDataE_26_port, 
                           y(25) => WriteDataE_25_port, y(24) => 
                           WriteDataE_24_port, y(23) => WriteDataE_23_port, 
                           y(22) => WriteDataE_22_port, y(21) => 
                           WriteDataE_21_port, y(20) => WriteDataE_20_port, 
                           y(19) => WriteDataE_19_port, y(18) => 
                           WriteDataE_18_port, y(17) => WriteDataE_17_port, 
                           y(16) => WriteDataE_16_port, y(15) => 
                           WriteDataE_15_port, y(14) => WriteDataE_14_port, 
                           y(13) => WriteDataE_13_port, y(12) => 
                           WriteDataE_12_port, y(11) => WriteDataE_11_port, 
                           y(10) => WriteDataE_10_port, y(9) => 
                           WriteDataE_9_port, y(8) => WriteDataE_8_port, y(7) 
                           => WriteDataE_7_port, y(6) => WriteDataE_6_port, 
                           y(5) => WriteDataE_5_port, y(4) => WriteDataE_4_port
                           , y(3) => WriteDataE_3_port, y(2) => 
                           WriteDataE_2_port, y(1) => WriteDataE_1_port, y(0) 
                           => WriteDataE_0_port);
   selSrcB : MUX21_N32_3 port map( a(31) => WriteDataE_31_port, a(30) => 
                           WriteDataE_30_port, a(29) => WriteDataE_29_port, 
                           a(28) => WriteDataE_28_port, a(27) => 
                           WriteDataE_27_port, a(26) => WriteDataE_26_port, 
                           a(25) => WriteDataE_25_port, a(24) => 
                           WriteDataE_24_port, a(23) => WriteDataE_23_port, 
                           a(22) => WriteDataE_22_port, a(21) => 
                           WriteDataE_21_port, a(20) => WriteDataE_20_port, 
                           a(19) => WriteDataE_19_port, a(18) => 
                           WriteDataE_18_port, a(17) => WriteDataE_17_port, 
                           a(16) => WriteDataE_16_port, a(15) => 
                           WriteDataE_15_port, a(14) => WriteDataE_14_port, 
                           a(13) => WriteDataE_13_port, a(12) => 
                           WriteDataE_12_port, a(11) => WriteDataE_11_port, 
                           a(10) => WriteDataE_10_port, a(9) => 
                           WriteDataE_9_port, a(8) => WriteDataE_8_port, a(7) 
                           => WriteDataE_7_port, a(6) => WriteDataE_6_port, 
                           a(5) => WriteDataE_5_port, a(4) => WriteDataE_4_port
                           , a(3) => WriteDataE_3_port, a(2) => 
                           WriteDataE_2_port, a(1) => WriteDataE_1_port, a(0) 
                           => WriteDataE_0_port, b(31) => SignImmE(31), b(30) 
                           => SignImmE(30), b(29) => SignImmE(29), b(28) => 
                           SignImmE(28), b(27) => SignImmE(27), b(26) => 
                           SignImmE(26), b(25) => SignImmE(25), b(24) => 
                           SignImmE(24), b(23) => SignImmE(23), b(22) => 
                           SignImmE(22), b(21) => SignImmE(21), b(20) => 
                           SignImmE(20), b(19) => SignImmE(19), b(18) => 
                           SignImmE(18), b(17) => SignImmE(17), b(16) => 
                           SignImmE(16), b(15) => SignImmE(15), b(14) => 
                           SignImmE(14), b(13) => SignImmE(13), b(12) => 
                           SignImmE(12), b(11) => SignImmE(11), b(10) => 
                           SignImmE(10), b(9) => SignImmE(9), b(8) => 
                           SignImmE(8), b(7) => SignImmE(7), b(6) => 
                           SignImmE(6), b(5) => SignImmE(5), b(4) => 
                           SignImmE(4), b(3) => SignImmE(3), b(2) => 
                           SignImmE(2), b(1) => SignImmE(1), b(0) => 
                           SignImmE(0), sel => ALUSrcE, y(31) => SrcBE_31_port,
                           y(30) => SrcBE_30_port, y(29) => SrcBE_29_port, 
                           y(28) => SrcBE_28_port, y(27) => SrcBE_27_port, 
                           y(26) => SrcBE_26_port, y(25) => SrcBE_25_port, 
                           y(24) => SrcBE_24_port, y(23) => SrcBE_23_port, 
                           y(22) => SrcBE_22_port, y(21) => SrcBE_21_port, 
                           y(20) => SrcBE_20_port, y(19) => SrcBE_19_port, 
                           y(18) => SrcBE_18_port, y(17) => SrcBE_17_port, 
                           y(16) => SrcBE_16_port, y(15) => SrcBE_15_port, 
                           y(14) => SrcBE_14_port, y(13) => SrcBE_13_port, 
                           y(12) => SrcBE_12_port, y(11) => SrcBE_11_port, 
                           y(10) => SrcBE_10_port, y(9) => SrcBE_9_port, y(8) 
                           => SrcBE_8_port, y(7) => SrcBE_7_port, y(6) => 
                           SrcBE_6_port, y(5) => SrcBE_5_port, y(4) => 
                           SrcBE_4_port, y(3) => SrcBE_3_port, y(2) => 
                           SrcBE_2_port, y(1) => SrcBE_1_port, y(0) => 
                           SrcBE_0_port);
   regAddr : MUX21_N5_1 port map( a(4) => RtE(4), a(3) => RtE(3), a(2) => 
                           RtE(2), a(1) => RtE(1), a(0) => RtE(0), b(4) => 
                           RdE(4), b(3) => RdE(3), b(2) => RdE(2), b(1) => 
                           RdE(1), b(0) => RdE(0), sel => RegDstE, y(4) => 
                           WriteRegE(4), y(3) => WriteRegE(3), y(2) => 
                           WriteRegE(2), y(1) => WriteRegE(1), y(0) => 
                           WriteRegE(0));
   ALUcomp : ALU_NBIT32 port map( en_alu => en_alu, op1(31) => SrcAE_31_port, 
                           op1(30) => SrcAE_30_port, op1(29) => SrcAE_29_port, 
                           op1(28) => SrcAE_28_port, op1(27) => SrcAE_27_port, 
                           op1(26) => SrcAE_26_port, op1(25) => SrcAE_25_port, 
                           op1(24) => SrcAE_24_port, op1(23) => SrcAE_23_port, 
                           op1(22) => SrcAE_22_port, op1(21) => SrcAE_21_port, 
                           op1(20) => SrcAE_20_port, op1(19) => SrcAE_19_port, 
                           op1(18) => SrcAE_18_port, op1(17) => SrcAE_17_port, 
                           op1(16) => SrcAE_16_port, op1(15) => SrcAE_15_port, 
                           op1(14) => SrcAE_14_port, op1(13) => SrcAE_13_port, 
                           op1(12) => SrcAE_12_port, op1(11) => SrcAE_11_port, 
                           op1(10) => SrcAE_10_port, op1(9) => SrcAE_9_port, 
                           op1(8) => SrcAE_8_port, op1(7) => SrcAE_7_port, 
                           op1(6) => SrcAE_6_port, op1(5) => SrcAE_5_port, 
                           op1(4) => SrcAE_4_port, op1(3) => SrcAE_3_port, 
                           op1(2) => SrcAE_2_port, op1(1) => SrcAE_1_port, 
                           op1(0) => SrcAE_0_port, op2(31) => SrcBE_31_port, 
                           op2(30) => SrcBE_30_port, op2(29) => SrcBE_29_port, 
                           op2(28) => SrcBE_28_port, op2(27) => SrcBE_27_port, 
                           op2(26) => SrcBE_26_port, op2(25) => SrcBE_25_port, 
                           op2(24) => SrcBE_24_port, op2(23) => SrcBE_23_port, 
                           op2(22) => SrcBE_22_port, op2(21) => SrcBE_21_port, 
                           op2(20) => SrcBE_20_port, op2(19) => SrcBE_19_port, 
                           op2(18) => SrcBE_18_port, op2(17) => SrcBE_17_port, 
                           op2(16) => SrcBE_16_port, op2(15) => SrcBE_15_port, 
                           op2(14) => SrcBE_14_port, op2(13) => SrcBE_13_port, 
                           op2(12) => SrcBE_12_port, op2(11) => SrcBE_11_port, 
                           op2(10) => SrcBE_10_port, op2(9) => SrcBE_9_port, 
                           op2(8) => SrcBE_8_port, op2(7) => SrcBE_7_port, 
                           op2(6) => SrcBE_6_port, op2(5) => SrcBE_5_port, 
                           op2(4) => SrcBE_4_port, op2(3) => SrcBE_3_port, 
                           op2(2) => SrcBE_2_port, op2(1) => SrcBE_1_port, 
                           op2(0) => SrcBE_0_port, sel(5) => ALUcontrolE(5), 
                           sel(4) => ALUcontrolE(4), sel(3) => ALUcontrolE(3), 
                           sel(2) => ALUcontrolE(2), sel(1) => ALUcontrolE(1), 
                           sel(0) => ALUcontrolE(0), result(31) => ALUoutE(31),
                           result(30) => ALUoutE(30), result(29) => ALUoutE(29)
                           , result(28) => ALUoutE(28), result(27) => 
                           ALUoutE(27), result(26) => ALUoutE(26), result(25) 
                           => ALUoutE(25), result(24) => ALUoutE(24), 
                           result(23) => ALUoutE(23), result(22) => ALUoutE(22)
                           , result(21) => ALUoutE(21), result(20) => 
                           ALUoutE(20), result(19) => ALUoutE(19), result(18) 
                           => ALUoutE(18), result(17) => ALUoutE(17), 
                           result(16) => ALUoutE(16), result(15) => ALUoutE(15)
                           , result(14) => ALUoutE(14), result(13) => 
                           ALUoutE(13), result(12) => ALUoutE(12), result(11) 
                           => ALUoutE(11), result(10) => ALUoutE(10), result(9)
                           => ALUoutE(9), result(8) => ALUoutE(8), result(7) =>
                           ALUoutE(7), result(6) => ALUoutE(6), result(5) => 
                           ALUoutE(5), result(4) => ALUoutE(4), result(3) => 
                           ALUoutE(3), result(2) => ALUoutE(2), result(1) => 
                           ALUoutE(1), result(0) => ALUoutE(0), CarryOut => 
                           n_1545, overflow => n_1546);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity Decode_wrapper is

   port( instrD, PcPlus4D : in std_logic_vector (31 downto 0);  select_ext, 
         ForwardAd, ForwardBD, clk, en, rst, RD1_EN, RD2_EN : in std_logic;  
         ALUOutM : in std_logic_vector (31 downto 0);  WriteRegW : in 
         std_logic_vector (4 downto 0);  ResultW : in std_logic_vector (31 
         downto 0);  CALL, RET, IsJal : in std_logic;  Comp_control : in 
         std_logic_vector (1 downto 0);  RegWriteW : in std_logic;  Memory_in :
         in std_logic_vector (31 downto 0);  Memory_out : out std_logic_vector 
         (31 downto 0);  FILL, SPILL : out std_logic;  RsD, RtD, RdE : out 
         std_logic_vector (4 downto 0);  SignImmD, PCBranchD : out 
         std_logic_vector (31 downto 0);  EqualD : out std_logic;  OP : out 
         std_logic_vector (5 downto 0);  FUNC : out std_logic_vector (10 downto
         0);  RD1, RD2 : out std_logic_vector (31 downto 0));

end Decode_wrapper;

architecture SYN_Behavioral of Decode_wrapper is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_addr
      port( y1, y2 : in std_logic_vector (31 downto 0);  comp_control : in 
            std_logic_vector (1 downto 0);  EqualD : out std_logic);
   end component;
   
   component MUX21_N32_4
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N32_5
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component window_rf_M4_N4_F4_NBIT32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  WR_ADD, RD1_ADD, 
            RD2_ADD : in std_logic_vector (4 downto 0);  FILL, SPILL : out 
            std_logic;  CALL, RET : in std_logic;  MEM_IN : in std_logic_vector
            (31 downto 0);  MEM_OUT : out std_logic_vector (31 downto 0);  
            DATAIN : in std_logic_vector (31 downto 0);  OUT1, OUT2 : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N5_0
      port( a, b : in std_logic_vector (4 downto 0);  sel : in std_logic;  y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component OR_GATE
      port( x, y : in std_logic;  z : out std_logic);
   end component;
   
   component MUX21_N32_6
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component adder_generic_nbit32
      port( a, b : in std_logic_vector (31 downto 0);  y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component sign_ext
      port( a : in std_logic_vector (31 downto 0);  s : in std_logic;  y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, SignImmD_31_port, SignImmD_30_port, SignImmD_29_port, 
      SignImmD_28_port, SignImmD_27_port, SignImmD_26_port, SignImmD_25_port, 
      SignImmD_24_port, SignImmD_23_port, SignImmD_22_port, SignImmD_21_port, 
      SignImmD_20_port, SignImmD_19_port, SignImmD_18_port, SignImmD_17_port, 
      SignImmD_16_port, SignImmD_15_port, SignImmD_14_port, SignImmD_13_port, 
      SignImmD_12_port, SignImmD_11_port, SignImmD_10_port, SignImmD_9_port, 
      SignImmD_8_port, SignImmD_7_port, SignImmD_6_port, SignImmD_5_port, 
      SignImmD_4_port, SignImmD_3_port, SignImmD_2_port, SignImmD_1_port, 
      SignImmD_0_port, RD1_31_port, RD1_30_port, RD1_29_port, RD1_28_port, 
      RD1_27_port, RD1_26_port, RD1_25_port, RD1_24_port, RD1_23_port, 
      RD1_22_port, RD1_21_port, RD1_20_port, RD1_19_port, RD1_18_port, 
      RD1_17_port, RD1_16_port, RD1_15_port, RD1_14_port, RD1_13_port, 
      RD1_12_port, RD1_11_port, RD1_10_port, RD1_9_port, RD1_8_port, RD1_7_port
      , RD1_6_port, RD1_5_port, RD1_4_port, RD1_3_port, RD1_2_port, RD1_1_port,
      RD1_0_port, RD2_31_port, RD2_30_port, RD2_29_port, RD2_28_port, 
      RD2_27_port, RD2_26_port, RD2_25_port, RD2_24_port, RD2_23_port, 
      RD2_22_port, RD2_21_port, RD2_20_port, RD2_19_port, RD2_18_port, 
      RD2_17_port, RD2_16_port, RD2_15_port, RD2_14_port, RD2_13_port, 
      RD2_12_port, RD2_11_port, RD2_10_port, RD2_9_port, RD2_8_port, RD2_7_port
      , RD2_6_port, RD2_5_port, RD2_4_port, RD2_3_port, RD2_2_port, RD2_1_port,
      RD2_0_port, ResultOrJal_31_port, ResultOrJal_30_port, ResultOrJal_29_port
      , ResultOrJal_28_port, ResultOrJal_27_port, ResultOrJal_26_port, 
      ResultOrJal_25_port, ResultOrJal_24_port, ResultOrJal_23_port, 
      ResultOrJal_22_port, ResultOrJal_21_port, ResultOrJal_20_port, 
      ResultOrJal_19_port, ResultOrJal_18_port, ResultOrJal_17_port, 
      ResultOrJal_16_port, ResultOrJal_15_port, ResultOrJal_14_port, 
      ResultOrJal_13_port, ResultOrJal_12_port, ResultOrJal_11_port, 
      ResultOrJal_10_port, ResultOrJal_9_port, ResultOrJal_8_port, 
      ResultOrJal_7_port, ResultOrJal_6_port, ResultOrJal_5_port, 
      ResultOrJal_4_port, ResultOrJal_3_port, ResultOrJal_2_port, 
      ResultOrJal_1_port, ResultOrJal_0_port, enable_for_W_RF, 
      Addr_or_R31_4_port, Addr_or_R31_3_port, Addr_or_R31_2_port, 
      Addr_or_R31_1_port, Addr_or_R31_0_port, RD1_rf_31_port, RD1_rf_30_port, 
      RD1_rf_29_port, RD1_rf_28_port, RD1_rf_27_port, RD1_rf_26_port, 
      RD1_rf_25_port, RD1_rf_24_port, RD1_rf_23_port, RD1_rf_22_port, 
      RD1_rf_21_port, RD1_rf_20_port, RD1_rf_19_port, RD1_rf_18_port, 
      RD1_rf_17_port, RD1_rf_16_port, RD1_rf_15_port, RD1_rf_14_port, 
      RD1_rf_13_port, RD1_rf_12_port, RD1_rf_11_port, RD1_rf_10_port, 
      RD1_rf_9_port, RD1_rf_8_port, RD1_rf_7_port, RD1_rf_6_port, RD1_rf_5_port
      , RD1_rf_4_port, RD1_rf_3_port, RD1_rf_2_port, RD1_rf_1_port, 
      RD1_rf_0_port, RD2_rf_31_port, RD2_rf_30_port, RD2_rf_29_port, 
      RD2_rf_28_port, RD2_rf_27_port, RD2_rf_26_port, RD2_rf_25_port, 
      RD2_rf_24_port, RD2_rf_23_port, RD2_rf_22_port, RD2_rf_21_port, 
      RD2_rf_20_port, RD2_rf_19_port, RD2_rf_18_port, RD2_rf_17_port, 
      RD2_rf_16_port, RD2_rf_15_port, RD2_rf_14_port, RD2_rf_13_port, 
      RD2_rf_12_port, RD2_rf_11_port, RD2_rf_10_port, RD2_rf_9_port, 
      RD2_rf_8_port, RD2_rf_7_port, RD2_rf_6_port, RD2_rf_5_port, RD2_rf_4_port
      , RD2_rf_3_port, RD2_rf_2_port, RD2_rf_1_port, RD2_rf_0_port, n1, n_1547 
      : std_logic;

begin
   RsD <= ( instrD(25), instrD(24), instrD(23), instrD(22), instrD(21) );
   RtD <= ( instrD(20), instrD(19), instrD(18), instrD(17), instrD(16) );
   RdE <= ( instrD(15), instrD(14), instrD(13), instrD(12), instrD(11) );
   SignImmD <= ( SignImmD_31_port, SignImmD_30_port, SignImmD_29_port, 
      SignImmD_28_port, SignImmD_27_port, SignImmD_26_port, SignImmD_25_port, 
      SignImmD_24_port, SignImmD_23_port, SignImmD_22_port, SignImmD_21_port, 
      SignImmD_20_port, SignImmD_19_port, SignImmD_18_port, SignImmD_17_port, 
      SignImmD_16_port, SignImmD_15_port, SignImmD_14_port, SignImmD_13_port, 
      SignImmD_12_port, SignImmD_11_port, SignImmD_10_port, SignImmD_9_port, 
      SignImmD_8_port, SignImmD_7_port, SignImmD_6_port, SignImmD_5_port, 
      SignImmD_4_port, SignImmD_3_port, SignImmD_2_port, SignImmD_1_port, 
      SignImmD_0_port );
   OP <= ( instrD(31), instrD(30), instrD(29), instrD(28), instrD(27), 
      instrD(26) );
   FUNC <= ( instrD(10), instrD(9), instrD(8), instrD(7), instrD(6), instrD(5),
      instrD(4), instrD(3), instrD(2), instrD(1), instrD(0) );
   RD1 <= ( RD1_31_port, RD1_30_port, RD1_29_port, RD1_28_port, RD1_27_port, 
      RD1_26_port, RD1_25_port, RD1_24_port, RD1_23_port, RD1_22_port, 
      RD1_21_port, RD1_20_port, RD1_19_port, RD1_18_port, RD1_17_port, 
      RD1_16_port, RD1_15_port, RD1_14_port, RD1_13_port, RD1_12_port, 
      RD1_11_port, RD1_10_port, RD1_9_port, RD1_8_port, RD1_7_port, RD1_6_port,
      RD1_5_port, RD1_4_port, RD1_3_port, RD1_2_port, RD1_1_port, RD1_0_port );
   RD2 <= ( RD2_31_port, RD2_30_port, RD2_29_port, RD2_28_port, RD2_27_port, 
      RD2_26_port, RD2_25_port, RD2_24_port, RD2_23_port, RD2_22_port, 
      RD2_21_port, RD2_20_port, RD2_19_port, RD2_18_port, RD2_17_port, 
      RD2_16_port, RD2_15_port, RD2_14_port, RD2_13_port, RD2_12_port, 
      RD2_11_port, RD2_10_port, RD2_9_port, RD2_8_port, RD2_7_port, RD2_6_port,
      RD2_5_port, RD2_4_port, RD2_3_port, RD2_2_port, RD2_1_port, RD2_0_port );
   
   X_Logic1_port <= '1';
   Sign_extended : sign_ext port map( a(31) => instrD(31), a(30) => instrD(30),
                           a(29) => instrD(29), a(28) => instrD(28), a(27) => 
                           instrD(27), a(26) => instrD(26), a(25) => instrD(25)
                           , a(24) => instrD(24), a(23) => instrD(23), a(22) =>
                           instrD(22), a(21) => instrD(21), a(20) => instrD(20)
                           , a(19) => instrD(19), a(18) => instrD(18), a(17) =>
                           instrD(17), a(16) => instrD(16), a(15) => instrD(15)
                           , a(14) => instrD(14), a(13) => instrD(13), a(12) =>
                           instrD(12), a(11) => instrD(11), a(10) => instrD(10)
                           , a(9) => instrD(9), a(8) => instrD(8), a(7) => 
                           instrD(7), a(6) => instrD(6), a(5) => instrD(5), 
                           a(4) => instrD(4), a(3) => instrD(3), a(2) => 
                           instrD(2), a(1) => instrD(1), a(0) => instrD(0), s 
                           => select_ext, y(31) => SignImmD_31_port, y(30) => 
                           SignImmD_30_port, y(29) => SignImmD_29_port, y(28) 
                           => SignImmD_28_port, y(27) => SignImmD_27_port, 
                           y(26) => SignImmD_26_port, y(25) => SignImmD_25_port
                           , y(24) => SignImmD_24_port, y(23) => 
                           SignImmD_23_port, y(22) => SignImmD_22_port, y(21) 
                           => SignImmD_21_port, y(20) => SignImmD_20_port, 
                           y(19) => SignImmD_19_port, y(18) => SignImmD_18_port
                           , y(17) => SignImmD_17_port, y(16) => 
                           SignImmD_16_port, y(15) => SignImmD_15_port, y(14) 
                           => SignImmD_14_port, y(13) => SignImmD_13_port, 
                           y(12) => SignImmD_12_port, y(11) => SignImmD_11_port
                           , y(10) => SignImmD_10_port, y(9) => SignImmD_9_port
                           , y(8) => SignImmD_8_port, y(7) => SignImmD_7_port, 
                           y(6) => SignImmD_6_port, y(5) => SignImmD_5_port, 
                           y(4) => SignImmD_4_port, y(3) => SignImmD_3_port, 
                           y(2) => SignImmD_2_port, y(1) => SignImmD_1_port, 
                           y(0) => SignImmD_0_port);
   adder : adder_generic_nbit32 port map( a(31) => SignImmD_31_port, a(30) => 
                           SignImmD_30_port, a(29) => SignImmD_29_port, a(28) 
                           => SignImmD_28_port, a(27) => SignImmD_27_port, 
                           a(26) => SignImmD_26_port, a(25) => SignImmD_25_port
                           , a(24) => SignImmD_24_port, a(23) => 
                           SignImmD_23_port, a(22) => SignImmD_22_port, a(21) 
                           => SignImmD_21_port, a(20) => SignImmD_20_port, 
                           a(19) => SignImmD_19_port, a(18) => SignImmD_18_port
                           , a(17) => SignImmD_17_port, a(16) => 
                           SignImmD_16_port, a(15) => SignImmD_15_port, a(14) 
                           => SignImmD_14_port, a(13) => SignImmD_13_port, 
                           a(12) => SignImmD_12_port, a(11) => SignImmD_11_port
                           , a(10) => SignImmD_10_port, a(9) => SignImmD_9_port
                           , a(8) => SignImmD_8_port, a(7) => SignImmD_7_port, 
                           a(6) => SignImmD_6_port, a(5) => SignImmD_5_port, 
                           a(4) => SignImmD_4_port, a(3) => SignImmD_3_port, 
                           a(2) => SignImmD_2_port, a(1) => SignImmD_1_port, 
                           a(0) => SignImmD_0_port, b(31) => PcPlus4D(31), 
                           b(30) => PcPlus4D(30), b(29) => PcPlus4D(29), b(28) 
                           => PcPlus4D(28), b(27) => PcPlus4D(27), b(26) => 
                           PcPlus4D(26), b(25) => PcPlus4D(25), b(24) => 
                           PcPlus4D(24), b(23) => PcPlus4D(23), b(22) => 
                           PcPlus4D(22), b(21) => PcPlus4D(21), b(20) => 
                           PcPlus4D(20), b(19) => PcPlus4D(19), b(18) => 
                           PcPlus4D(18), b(17) => PcPlus4D(17), b(16) => 
                           PcPlus4D(16), b(15) => PcPlus4D(15), b(14) => 
                           PcPlus4D(14), b(13) => PcPlus4D(13), b(12) => 
                           PcPlus4D(12), b(11) => PcPlus4D(11), b(10) => 
                           PcPlus4D(10), b(9) => PcPlus4D(9), b(8) => 
                           PcPlus4D(8), b(7) => PcPlus4D(7), b(6) => 
                           PcPlus4D(6), b(5) => PcPlus4D(5), b(4) => 
                           PcPlus4D(4), b(3) => PcPlus4D(3), b(2) => 
                           PcPlus4D(2), b(1) => PcPlus4D(1), b(0) => 
                           PcPlus4D(0), y(31) => PCBranchD(31), y(30) => 
                           PCBranchD(30), y(29) => PCBranchD(29), y(28) => 
                           PCBranchD(28), y(27) => PCBranchD(27), y(26) => 
                           PCBranchD(26), y(25) => PCBranchD(25), y(24) => 
                           PCBranchD(24), y(23) => PCBranchD(23), y(22) => 
                           PCBranchD(22), y(21) => PCBranchD(21), y(20) => 
                           PCBranchD(20), y(19) => PCBranchD(19), y(18) => 
                           PCBranchD(18), y(17) => PCBranchD(17), y(16) => 
                           PCBranchD(16), y(15) => PCBranchD(15), y(14) => 
                           PCBranchD(14), y(13) => PCBranchD(13), y(12) => 
                           PCBranchD(12), y(11) => PCBranchD(11), y(10) => 
                           PCBranchD(10), y(9) => PCBranchD(9), y(8) => 
                           PCBranchD(8), y(7) => PCBranchD(7), y(6) => 
                           PCBranchD(6), y(5) => PCBranchD(5), y(4) => 
                           PCBranchD(4), y(3) => PCBranchD(3), y(2) => 
                           PCBranchD(2), y(1) => PCBranchD(1), y(0) => 
                           PCBranchD(0));
   MUX3 : MUX21_N32_6 port map( a(31) => ResultW(31), a(30) => ResultW(30), 
                           a(29) => ResultW(29), a(28) => ResultW(28), a(27) =>
                           ResultW(27), a(26) => ResultW(26), a(25) => 
                           ResultW(25), a(24) => ResultW(24), a(23) => 
                           ResultW(23), a(22) => ResultW(22), a(21) => 
                           ResultW(21), a(20) => ResultW(20), a(19) => 
                           ResultW(19), a(18) => ResultW(18), a(17) => 
                           ResultW(17), a(16) => ResultW(16), a(15) => 
                           ResultW(15), a(14) => ResultW(14), a(13) => 
                           ResultW(13), a(12) => ResultW(12), a(11) => 
                           ResultW(11), a(10) => ResultW(10), a(9) => 
                           ResultW(9), a(8) => ResultW(8), a(7) => ResultW(7), 
                           a(6) => ResultW(6), a(5) => ResultW(5), a(4) => 
                           ResultW(4), a(3) => ResultW(3), a(2) => ResultW(2), 
                           a(1) => ResultW(1), a(0) => ResultW(0), b(31) => 
                           PcPlus4D(31), b(30) => PcPlus4D(30), b(29) => 
                           PcPlus4D(29), b(28) => PcPlus4D(28), b(27) => 
                           PcPlus4D(27), b(26) => PcPlus4D(26), b(25) => 
                           PcPlus4D(25), b(24) => PcPlus4D(24), b(23) => 
                           PcPlus4D(23), b(22) => PcPlus4D(22), b(21) => 
                           PcPlus4D(21), b(20) => PcPlus4D(20), b(19) => 
                           PcPlus4D(19), b(18) => PcPlus4D(18), b(17) => 
                           PcPlus4D(17), b(16) => PcPlus4D(16), b(15) => 
                           PcPlus4D(15), b(14) => PcPlus4D(14), b(13) => 
                           PcPlus4D(13), b(12) => PcPlus4D(12), b(11) => 
                           PcPlus4D(11), b(10) => PcPlus4D(10), b(9) => 
                           PcPlus4D(9), b(8) => PcPlus4D(8), b(7) => 
                           PcPlus4D(7), b(6) => PcPlus4D(6), b(5) => 
                           PcPlus4D(5), b(4) => PcPlus4D(4), b(3) => 
                           PcPlus4D(3), b(2) => PcPlus4D(2), b(1) => 
                           PcPlus4D(1), b(0) => PcPlus4D(0), sel => IsJal, 
                           y(31) => ResultOrJal_31_port, y(30) => 
                           ResultOrJal_30_port, y(29) => ResultOrJal_29_port, 
                           y(28) => ResultOrJal_28_port, y(27) => 
                           ResultOrJal_27_port, y(26) => ResultOrJal_26_port, 
                           y(25) => ResultOrJal_25_port, y(24) => 
                           ResultOrJal_24_port, y(23) => ResultOrJal_23_port, 
                           y(22) => ResultOrJal_22_port, y(21) => 
                           ResultOrJal_21_port, y(20) => ResultOrJal_20_port, 
                           y(19) => ResultOrJal_19_port, y(18) => 
                           ResultOrJal_18_port, y(17) => ResultOrJal_17_port, 
                           y(16) => ResultOrJal_16_port, y(15) => 
                           ResultOrJal_15_port, y(14) => ResultOrJal_14_port, 
                           y(13) => ResultOrJal_13_port, y(12) => 
                           ResultOrJal_12_port, y(11) => ResultOrJal_11_port, 
                           y(10) => ResultOrJal_10_port, y(9) => 
                           ResultOrJal_9_port, y(8) => ResultOrJal_8_port, y(7)
                           => ResultOrJal_7_port, y(6) => ResultOrJal_6_port, 
                           y(5) => ResultOrJal_5_port, y(4) => 
                           ResultOrJal_4_port, y(3) => ResultOrJal_3_port, y(2)
                           => ResultOrJal_2_port, y(1) => ResultOrJal_1_port, 
                           y(0) => ResultOrJal_0_port);
   OR1 : OR_GATE port map( x => IsJal, y => RegWriteW, z => enable_for_W_RF);
   MUX4 : MUX21_N5_0 port map( a(4) => WriteRegW(4), a(3) => WriteRegW(3), a(2)
                           => WriteRegW(2), a(1) => WriteRegW(1), a(0) => 
                           WriteRegW(0), b(4) => X_Logic1_port, b(3) => 
                           X_Logic1_port, b(2) => X_Logic1_port, b(1) => 
                           X_Logic1_port, b(0) => X_Logic1_port, sel => IsJal, 
                           y(4) => Addr_or_R31_4_port, y(3) => 
                           Addr_or_R31_3_port, y(2) => Addr_or_R31_2_port, y(1)
                           => Addr_or_R31_1_port, y(0) => Addr_or_R31_0_port);
   RF : window_rf_M4_N4_F4_NBIT32 port map( CLK => n1, RESET => rst, ENABLE => 
                           en, RD1 => RD1_EN, RD2 => RD2_EN, WR => 
                           enable_for_W_RF, WR_ADD(4) => Addr_or_R31_4_port, 
                           WR_ADD(3) => Addr_or_R31_3_port, WR_ADD(2) => 
                           Addr_or_R31_2_port, WR_ADD(1) => Addr_or_R31_1_port,
                           WR_ADD(0) => Addr_or_R31_0_port, RD1_ADD(4) => 
                           instrD(25), RD1_ADD(3) => instrD(24), RD1_ADD(2) => 
                           instrD(23), RD1_ADD(1) => instrD(22), RD1_ADD(0) => 
                           instrD(21), RD2_ADD(4) => instrD(20), RD2_ADD(3) => 
                           instrD(19), RD2_ADD(2) => instrD(18), RD2_ADD(1) => 
                           instrD(17), RD2_ADD(0) => instrD(16), FILL => FILL, 
                           SPILL => n_1547, CALL => CALL, RET => RET, 
                           MEM_IN(31) => Memory_in(31), MEM_IN(30) => 
                           Memory_in(30), MEM_IN(29) => Memory_in(29), 
                           MEM_IN(28) => Memory_in(28), MEM_IN(27) => 
                           Memory_in(27), MEM_IN(26) => Memory_in(26), 
                           MEM_IN(25) => Memory_in(25), MEM_IN(24) => 
                           Memory_in(24), MEM_IN(23) => Memory_in(23), 
                           MEM_IN(22) => Memory_in(22), MEM_IN(21) => 
                           Memory_in(21), MEM_IN(20) => Memory_in(20), 
                           MEM_IN(19) => Memory_in(19), MEM_IN(18) => 
                           Memory_in(18), MEM_IN(17) => Memory_in(17), 
                           MEM_IN(16) => Memory_in(16), MEM_IN(15) => 
                           Memory_in(15), MEM_IN(14) => Memory_in(14), 
                           MEM_IN(13) => Memory_in(13), MEM_IN(12) => 
                           Memory_in(12), MEM_IN(11) => Memory_in(11), 
                           MEM_IN(10) => Memory_in(10), MEM_IN(9) => 
                           Memory_in(9), MEM_IN(8) => Memory_in(8), MEM_IN(7) 
                           => Memory_in(7), MEM_IN(6) => Memory_in(6), 
                           MEM_IN(5) => Memory_in(5), MEM_IN(4) => Memory_in(4)
                           , MEM_IN(3) => Memory_in(3), MEM_IN(2) => 
                           Memory_in(2), MEM_IN(1) => Memory_in(1), MEM_IN(0) 
                           => Memory_in(0), MEM_OUT(31) => Memory_out(31), 
                           MEM_OUT(30) => Memory_out(30), MEM_OUT(29) => 
                           Memory_out(29), MEM_OUT(28) => Memory_out(28), 
                           MEM_OUT(27) => Memory_out(27), MEM_OUT(26) => 
                           Memory_out(26), MEM_OUT(25) => Memory_out(25), 
                           MEM_OUT(24) => Memory_out(24), MEM_OUT(23) => 
                           Memory_out(23), MEM_OUT(22) => Memory_out(22), 
                           MEM_OUT(21) => Memory_out(21), MEM_OUT(20) => 
                           Memory_out(20), MEM_OUT(19) => Memory_out(19), 
                           MEM_OUT(18) => Memory_out(18), MEM_OUT(17) => 
                           Memory_out(17), MEM_OUT(16) => Memory_out(16), 
                           MEM_OUT(15) => Memory_out(15), MEM_OUT(14) => 
                           Memory_out(14), MEM_OUT(13) => Memory_out(13), 
                           MEM_OUT(12) => Memory_out(12), MEM_OUT(11) => 
                           Memory_out(11), MEM_OUT(10) => Memory_out(10), 
                           MEM_OUT(9) => Memory_out(9), MEM_OUT(8) => 
                           Memory_out(8), MEM_OUT(7) => Memory_out(7), 
                           MEM_OUT(6) => Memory_out(6), MEM_OUT(5) => 
                           Memory_out(5), MEM_OUT(4) => Memory_out(4), 
                           MEM_OUT(3) => Memory_out(3), MEM_OUT(2) => 
                           Memory_out(2), MEM_OUT(1) => Memory_out(1), 
                           MEM_OUT(0) => Memory_out(0), DATAIN(31) => 
                           ResultOrJal_31_port, DATAIN(30) => 
                           ResultOrJal_30_port, DATAIN(29) => 
                           ResultOrJal_29_port, DATAIN(28) => 
                           ResultOrJal_28_port, DATAIN(27) => 
                           ResultOrJal_27_port, DATAIN(26) => 
                           ResultOrJal_26_port, DATAIN(25) => 
                           ResultOrJal_25_port, DATAIN(24) => 
                           ResultOrJal_24_port, DATAIN(23) => 
                           ResultOrJal_23_port, DATAIN(22) => 
                           ResultOrJal_22_port, DATAIN(21) => 
                           ResultOrJal_21_port, DATAIN(20) => 
                           ResultOrJal_20_port, DATAIN(19) => 
                           ResultOrJal_19_port, DATAIN(18) => 
                           ResultOrJal_18_port, DATAIN(17) => 
                           ResultOrJal_17_port, DATAIN(16) => 
                           ResultOrJal_16_port, DATAIN(15) => 
                           ResultOrJal_15_port, DATAIN(14) => 
                           ResultOrJal_14_port, DATAIN(13) => 
                           ResultOrJal_13_port, DATAIN(12) => 
                           ResultOrJal_12_port, DATAIN(11) => 
                           ResultOrJal_11_port, DATAIN(10) => 
                           ResultOrJal_10_port, DATAIN(9) => ResultOrJal_9_port
                           , DATAIN(8) => ResultOrJal_8_port, DATAIN(7) => 
                           ResultOrJal_7_port, DATAIN(6) => ResultOrJal_6_port,
                           DATAIN(5) => ResultOrJal_5_port, DATAIN(4) => 
                           ResultOrJal_4_port, DATAIN(3) => ResultOrJal_3_port,
                           DATAIN(2) => ResultOrJal_2_port, DATAIN(1) => 
                           ResultOrJal_1_port, DATAIN(0) => ResultOrJal_0_port,
                           OUT1(31) => RD1_rf_31_port, OUT1(30) => 
                           RD1_rf_30_port, OUT1(29) => RD1_rf_29_port, OUT1(28)
                           => RD1_rf_28_port, OUT1(27) => RD1_rf_27_port, 
                           OUT1(26) => RD1_rf_26_port, OUT1(25) => 
                           RD1_rf_25_port, OUT1(24) => RD1_rf_24_port, OUT1(23)
                           => RD1_rf_23_port, OUT1(22) => RD1_rf_22_port, 
                           OUT1(21) => RD1_rf_21_port, OUT1(20) => 
                           RD1_rf_20_port, OUT1(19) => RD1_rf_19_port, OUT1(18)
                           => RD1_rf_18_port, OUT1(17) => RD1_rf_17_port, 
                           OUT1(16) => RD1_rf_16_port, OUT1(15) => 
                           RD1_rf_15_port, OUT1(14) => RD1_rf_14_port, OUT1(13)
                           => RD1_rf_13_port, OUT1(12) => RD1_rf_12_port, 
                           OUT1(11) => RD1_rf_11_port, OUT1(10) => 
                           RD1_rf_10_port, OUT1(9) => RD1_rf_9_port, OUT1(8) =>
                           RD1_rf_8_port, OUT1(7) => RD1_rf_7_port, OUT1(6) => 
                           RD1_rf_6_port, OUT1(5) => RD1_rf_5_port, OUT1(4) => 
                           RD1_rf_4_port, OUT1(3) => RD1_rf_3_port, OUT1(2) => 
                           RD1_rf_2_port, OUT1(1) => RD1_rf_1_port, OUT1(0) => 
                           RD1_rf_0_port, OUT2(31) => RD2_rf_31_port, OUT2(30) 
                           => RD2_rf_30_port, OUT2(29) => RD2_rf_29_port, 
                           OUT2(28) => RD2_rf_28_port, OUT2(27) => 
                           RD2_rf_27_port, OUT2(26) => RD2_rf_26_port, OUT2(25)
                           => RD2_rf_25_port, OUT2(24) => RD2_rf_24_port, 
                           OUT2(23) => RD2_rf_23_port, OUT2(22) => 
                           RD2_rf_22_port, OUT2(21) => RD2_rf_21_port, OUT2(20)
                           => RD2_rf_20_port, OUT2(19) => RD2_rf_19_port, 
                           OUT2(18) => RD2_rf_18_port, OUT2(17) => 
                           RD2_rf_17_port, OUT2(16) => RD2_rf_16_port, OUT2(15)
                           => RD2_rf_15_port, OUT2(14) => RD2_rf_14_port, 
                           OUT2(13) => RD2_rf_13_port, OUT2(12) => 
                           RD2_rf_12_port, OUT2(11) => RD2_rf_11_port, OUT2(10)
                           => RD2_rf_10_port, OUT2(9) => RD2_rf_9_port, OUT2(8)
                           => RD2_rf_8_port, OUT2(7) => RD2_rf_7_port, OUT2(6) 
                           => RD2_rf_6_port, OUT2(5) => RD2_rf_5_port, OUT2(4) 
                           => RD2_rf_4_port, OUT2(3) => RD2_rf_3_port, OUT2(2) 
                           => RD2_rf_2_port, OUT2(1) => RD2_rf_1_port, OUT2(0) 
                           => RD2_rf_0_port);
   MUX1 : MUX21_N32_5 port map( a(31) => RD1_rf_31_port, a(30) => 
                           RD1_rf_30_port, a(29) => RD1_rf_29_port, a(28) => 
                           RD1_rf_28_port, a(27) => RD1_rf_27_port, a(26) => 
                           RD1_rf_26_port, a(25) => RD1_rf_25_port, a(24) => 
                           RD1_rf_24_port, a(23) => RD1_rf_23_port, a(22) => 
                           RD1_rf_22_port, a(21) => RD1_rf_21_port, a(20) => 
                           RD1_rf_20_port, a(19) => RD1_rf_19_port, a(18) => 
                           RD1_rf_18_port, a(17) => RD1_rf_17_port, a(16) => 
                           RD1_rf_16_port, a(15) => RD1_rf_15_port, a(14) => 
                           RD1_rf_14_port, a(13) => RD1_rf_13_port, a(12) => 
                           RD1_rf_12_port, a(11) => RD1_rf_11_port, a(10) => 
                           RD1_rf_10_port, a(9) => RD1_rf_9_port, a(8) => 
                           RD1_rf_8_port, a(7) => RD1_rf_7_port, a(6) => 
                           RD1_rf_6_port, a(5) => RD1_rf_5_port, a(4) => 
                           RD1_rf_4_port, a(3) => RD1_rf_3_port, a(2) => 
                           RD1_rf_2_port, a(1) => RD1_rf_1_port, a(0) => 
                           RD1_rf_0_port, b(31) => ALUOutM(31), b(30) => 
                           ALUOutM(30), b(29) => ALUOutM(29), b(28) => 
                           ALUOutM(28), b(27) => ALUOutM(27), b(26) => 
                           ALUOutM(26), b(25) => ALUOutM(25), b(24) => 
                           ALUOutM(24), b(23) => ALUOutM(23), b(22) => 
                           ALUOutM(22), b(21) => ALUOutM(21), b(20) => 
                           ALUOutM(20), b(19) => ALUOutM(19), b(18) => 
                           ALUOutM(18), b(17) => ALUOutM(17), b(16) => 
                           ALUOutM(16), b(15) => ALUOutM(15), b(14) => 
                           ALUOutM(14), b(13) => ALUOutM(13), b(12) => 
                           ALUOutM(12), b(11) => ALUOutM(11), b(10) => 
                           ALUOutM(10), b(9) => ALUOutM(9), b(8) => ALUOutM(8),
                           b(7) => ALUOutM(7), b(6) => ALUOutM(6), b(5) => 
                           ALUOutM(5), b(4) => ALUOutM(4), b(3) => ALUOutM(3), 
                           b(2) => ALUOutM(2), b(1) => ALUOutM(1), b(0) => 
                           ALUOutM(0), sel => ForwardAd, y(31) => RD1_31_port, 
                           y(30) => RD1_30_port, y(29) => RD1_29_port, y(28) =>
                           RD1_28_port, y(27) => RD1_27_port, y(26) => 
                           RD1_26_port, y(25) => RD1_25_port, y(24) => 
                           RD1_24_port, y(23) => RD1_23_port, y(22) => 
                           RD1_22_port, y(21) => RD1_21_port, y(20) => 
                           RD1_20_port, y(19) => RD1_19_port, y(18) => 
                           RD1_18_port, y(17) => RD1_17_port, y(16) => 
                           RD1_16_port, y(15) => RD1_15_port, y(14) => 
                           RD1_14_port, y(13) => RD1_13_port, y(12) => 
                           RD1_12_port, y(11) => RD1_11_port, y(10) => 
                           RD1_10_port, y(9) => RD1_9_port, y(8) => RD1_8_port,
                           y(7) => RD1_7_port, y(6) => RD1_6_port, y(5) => 
                           RD1_5_port, y(4) => RD1_4_port, y(3) => RD1_3_port, 
                           y(2) => RD1_2_port, y(1) => RD1_1_port, y(0) => 
                           RD1_0_port);
   MUX2 : MUX21_N32_4 port map( a(31) => RD2_rf_31_port, a(30) => 
                           RD2_rf_30_port, a(29) => RD2_rf_29_port, a(28) => 
                           RD2_rf_28_port, a(27) => RD2_rf_27_port, a(26) => 
                           RD2_rf_26_port, a(25) => RD2_rf_25_port, a(24) => 
                           RD2_rf_24_port, a(23) => RD2_rf_23_port, a(22) => 
                           RD2_rf_22_port, a(21) => RD2_rf_21_port, a(20) => 
                           RD2_rf_20_port, a(19) => RD2_rf_19_port, a(18) => 
                           RD2_rf_18_port, a(17) => RD2_rf_17_port, a(16) => 
                           RD2_rf_16_port, a(15) => RD2_rf_15_port, a(14) => 
                           RD2_rf_14_port, a(13) => RD2_rf_13_port, a(12) => 
                           RD2_rf_12_port, a(11) => RD2_rf_11_port, a(10) => 
                           RD2_rf_10_port, a(9) => RD2_rf_9_port, a(8) => 
                           RD2_rf_8_port, a(7) => RD2_rf_7_port, a(6) => 
                           RD2_rf_6_port, a(5) => RD2_rf_5_port, a(4) => 
                           RD2_rf_4_port, a(3) => RD2_rf_3_port, a(2) => 
                           RD2_rf_2_port, a(1) => RD2_rf_1_port, a(0) => 
                           RD2_rf_0_port, b(31) => ALUOutM(31), b(30) => 
                           ALUOutM(30), b(29) => ALUOutM(29), b(28) => 
                           ALUOutM(28), b(27) => ALUOutM(27), b(26) => 
                           ALUOutM(26), b(25) => ALUOutM(25), b(24) => 
                           ALUOutM(24), b(23) => ALUOutM(23), b(22) => 
                           ALUOutM(22), b(21) => ALUOutM(21), b(20) => 
                           ALUOutM(20), b(19) => ALUOutM(19), b(18) => 
                           ALUOutM(18), b(17) => ALUOutM(17), b(16) => 
                           ALUOutM(16), b(15) => ALUOutM(15), b(14) => 
                           ALUOutM(14), b(13) => ALUOutM(13), b(12) => 
                           ALUOutM(12), b(11) => ALUOutM(11), b(10) => 
                           ALUOutM(10), b(9) => ALUOutM(9), b(8) => ALUOutM(8),
                           b(7) => ALUOutM(7), b(6) => ALUOutM(6), b(5) => 
                           ALUOutM(5), b(4) => ALUOutM(4), b(3) => ALUOutM(3), 
                           b(2) => ALUOutM(2), b(1) => ALUOutM(1), b(0) => 
                           ALUOutM(0), sel => ForwardBD, y(31) => RD2_31_port, 
                           y(30) => RD2_30_port, y(29) => RD2_29_port, y(28) =>
                           RD2_28_port, y(27) => RD2_27_port, y(26) => 
                           RD2_26_port, y(25) => RD2_25_port, y(24) => 
                           RD2_24_port, y(23) => RD2_23_port, y(22) => 
                           RD2_22_port, y(21) => RD2_21_port, y(20) => 
                           RD2_20_port, y(19) => RD2_19_port, y(18) => 
                           RD2_18_port, y(17) => RD2_17_port, y(16) => 
                           RD2_16_port, y(15) => RD2_15_port, y(14) => 
                           RD2_14_port, y(13) => RD2_13_port, y(12) => 
                           RD2_12_port, y(11) => RD2_11_port, y(10) => 
                           RD2_10_port, y(9) => RD2_9_port, y(8) => RD2_8_port,
                           y(7) => RD2_7_port, y(6) => RD2_6_port, y(5) => 
                           RD2_5_port, y(4) => RD2_4_port, y(3) => RD2_3_port, 
                           y(2) => RD2_2_port, y(1) => RD2_1_port, y(0) => 
                           RD2_0_port);
   Comparator : comparator_addr port map( y1(31) => RD1_31_port, y1(30) => 
                           RD1_30_port, y1(29) => RD1_29_port, y1(28) => 
                           RD1_28_port, y1(27) => RD1_27_port, y1(26) => 
                           RD1_26_port, y1(25) => RD1_25_port, y1(24) => 
                           RD1_24_port, y1(23) => RD1_23_port, y1(22) => 
                           RD1_22_port, y1(21) => RD1_21_port, y1(20) => 
                           RD1_20_port, y1(19) => RD1_19_port, y1(18) => 
                           RD1_18_port, y1(17) => RD1_17_port, y1(16) => 
                           RD1_16_port, y1(15) => RD1_15_port, y1(14) => 
                           RD1_14_port, y1(13) => RD1_13_port, y1(12) => 
                           RD1_12_port, y1(11) => RD1_11_port, y1(10) => 
                           RD1_10_port, y1(9) => RD1_9_port, y1(8) => 
                           RD1_8_port, y1(7) => RD1_7_port, y1(6) => RD1_6_port
                           , y1(5) => RD1_5_port, y1(4) => RD1_4_port, y1(3) =>
                           RD1_3_port, y1(2) => RD1_2_port, y1(1) => RD1_1_port
                           , y1(0) => RD1_0_port, y2(31) => RD2_31_port, y2(30)
                           => RD2_30_port, y2(29) => RD2_29_port, y2(28) => 
                           RD2_28_port, y2(27) => RD2_27_port, y2(26) => 
                           RD2_26_port, y2(25) => RD2_25_port, y2(24) => 
                           RD2_24_port, y2(23) => RD2_23_port, y2(22) => 
                           RD2_22_port, y2(21) => RD2_21_port, y2(20) => 
                           RD2_20_port, y2(19) => RD2_19_port, y2(18) => 
                           RD2_18_port, y2(17) => RD2_17_port, y2(16) => 
                           RD2_16_port, y2(15) => RD2_15_port, y2(14) => 
                           RD2_14_port, y2(13) => RD2_13_port, y2(12) => 
                           RD2_12_port, y2(11) => RD2_11_port, y2(10) => 
                           RD2_10_port, y2(9) => RD2_9_port, y2(8) => 
                           RD2_8_port, y2(7) => RD2_7_port, y2(6) => RD2_6_port
                           , y2(5) => RD2_5_port, y2(4) => RD2_4_port, y2(3) =>
                           RD2_3_port, y2(2) => RD2_2_port, y2(1) => RD2_1_port
                           , y2(0) => RD2_0_port, comp_control(1) => 
                           Comp_control(1), comp_control(0) => Comp_control(0),
                           EqualD => EqualD);
   U2 : INV_X1 port map( A => clk, ZN => n1);
   SPILL <= '0';

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity fetch_stage_wrapper_nbit32_nwords64 is

   port( PCBranchD : in std_logic_vector (31 downto 0);  PCPlus4F, InstrD, 
         address_to_iram : out std_logic_vector (31 downto 0);  iram_to_dlx : 
         in std_logic_vector (31 downto 0);  PCSrcD, StallF, clk, rst : in 
         std_logic);

end fetch_stage_wrapper_nbit32_nwords64;

architecture SYN_structural of fetch_stage_wrapper_nbit32_nwords64 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component adder_genericu_nbit32
      port( a, b : in std_logic_vector (31 downto 0);  y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component register_generic_nbit32
      port( d : in std_logic_vector (31 downto 0);  q : out std_logic_vector 
            (31 downto 0);  clk, reset, en : in std_logic);
   end component;
   
   component MUX21_N32_0
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, PCPlus4F_31_port, PCPlus4F_30_port, 
      PCPlus4F_29_port, PCPlus4F_28_port, PCPlus4F_27_port, PCPlus4F_26_port, 
      PCPlus4F_25_port, PCPlus4F_24_port, PCPlus4F_23_port, PCPlus4F_22_port, 
      PCPlus4F_21_port, PCPlus4F_20_port, PCPlus4F_19_port, PCPlus4F_18_port, 
      PCPlus4F_17_port, PCPlus4F_16_port, PCPlus4F_15_port, PCPlus4F_14_port, 
      PCPlus4F_13_port, PCPlus4F_12_port, PCPlus4F_11_port, PCPlus4F_10_port, 
      PCPlus4F_9_port, PCPlus4F_8_port, PCPlus4F_7_port, PCPlus4F_6_port, 
      PCPlus4F_5_port, PCPlus4F_4_port, PCPlus4F_3_port, PCPlus4F_2_port, 
      PCPlus4F_1_port, PCPlus4F_0_port, address_to_iram_31_port, 
      address_to_iram_30_port, address_to_iram_29_port, address_to_iram_28_port
      , address_to_iram_27_port, address_to_iram_26_port, 
      address_to_iram_25_port, address_to_iram_24_port, address_to_iram_23_port
      , address_to_iram_22_port, address_to_iram_21_port, 
      address_to_iram_20_port, address_to_iram_19_port, address_to_iram_18_port
      , address_to_iram_17_port, address_to_iram_16_port, 
      address_to_iram_15_port, address_to_iram_14_port, address_to_iram_13_port
      , address_to_iram_12_port, address_to_iram_11_port, 
      address_to_iram_10_port, address_to_iram_9_port, address_to_iram_8_port, 
      address_to_iram_7_port, address_to_iram_6_port, address_to_iram_5_port, 
      address_to_iram_4_port, address_to_iram_3_port, address_to_iram_2_port, 
      address_to_iram_1_port, address_to_iram_0_port, PC_31_port, PC_30_port, 
      PC_29_port, PC_28_port, PC_27_port, PC_26_port, PC_25_port, PC_24_port, 
      PC_23_port, PC_22_port, PC_21_port, PC_20_port, PC_19_port, PC_18_port, 
      PC_17_port, PC_16_port, PC_15_port, PC_14_port, PC_13_port, PC_12_port, 
      PC_11_port, PC_10_port, PC_9_port, PC_8_port, PC_7_port, PC_6_port, 
      PC_5_port, PC_4_port, PC_3_port, PC_2_port, PC_1_port, PC_0_port, n1 : 
      std_logic;

begin
   PCPlus4F <= ( PCPlus4F_31_port, PCPlus4F_30_port, PCPlus4F_29_port, 
      PCPlus4F_28_port, PCPlus4F_27_port, PCPlus4F_26_port, PCPlus4F_25_port, 
      PCPlus4F_24_port, PCPlus4F_23_port, PCPlus4F_22_port, PCPlus4F_21_port, 
      PCPlus4F_20_port, PCPlus4F_19_port, PCPlus4F_18_port, PCPlus4F_17_port, 
      PCPlus4F_16_port, PCPlus4F_15_port, PCPlus4F_14_port, PCPlus4F_13_port, 
      PCPlus4F_12_port, PCPlus4F_11_port, PCPlus4F_10_port, PCPlus4F_9_port, 
      PCPlus4F_8_port, PCPlus4F_7_port, PCPlus4F_6_port, PCPlus4F_5_port, 
      PCPlus4F_4_port, PCPlus4F_3_port, PCPlus4F_2_port, PCPlus4F_1_port, 
      PCPlus4F_0_port );
   InstrD <= ( iram_to_dlx(31), iram_to_dlx(30), iram_to_dlx(29), 
      iram_to_dlx(28), iram_to_dlx(27), iram_to_dlx(26), iram_to_dlx(25), 
      iram_to_dlx(24), iram_to_dlx(23), iram_to_dlx(22), iram_to_dlx(21), 
      iram_to_dlx(20), iram_to_dlx(19), iram_to_dlx(18), iram_to_dlx(17), 
      iram_to_dlx(16), iram_to_dlx(15), iram_to_dlx(14), iram_to_dlx(13), 
      iram_to_dlx(12), iram_to_dlx(11), iram_to_dlx(10), iram_to_dlx(9), 
      iram_to_dlx(8), iram_to_dlx(7), iram_to_dlx(6), iram_to_dlx(5), 
      iram_to_dlx(4), iram_to_dlx(3), iram_to_dlx(2), iram_to_dlx(1), 
      iram_to_dlx(0) );
   address_to_iram <= ( address_to_iram_31_port, address_to_iram_30_port, 
      address_to_iram_29_port, address_to_iram_28_port, address_to_iram_27_port
      , address_to_iram_26_port, address_to_iram_25_port, 
      address_to_iram_24_port, address_to_iram_23_port, address_to_iram_22_port
      , address_to_iram_21_port, address_to_iram_20_port, 
      address_to_iram_19_port, address_to_iram_18_port, address_to_iram_17_port
      , address_to_iram_16_port, address_to_iram_15_port, 
      address_to_iram_14_port, address_to_iram_13_port, address_to_iram_12_port
      , address_to_iram_11_port, address_to_iram_10_port, 
      address_to_iram_9_port, address_to_iram_8_port, address_to_iram_7_port, 
      address_to_iram_6_port, address_to_iram_5_port, address_to_iram_4_port, 
      address_to_iram_3_port, address_to_iram_2_port, address_to_iram_1_port, 
      address_to_iram_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   pc_mux : MUX21_N32_0 port map( a(31) => PCPlus4F_31_port, a(30) => 
                           PCPlus4F_30_port, a(29) => PCPlus4F_29_port, a(28) 
                           => PCPlus4F_28_port, a(27) => PCPlus4F_27_port, 
                           a(26) => PCPlus4F_26_port, a(25) => PCPlus4F_25_port
                           , a(24) => PCPlus4F_24_port, a(23) => 
                           PCPlus4F_23_port, a(22) => PCPlus4F_22_port, a(21) 
                           => PCPlus4F_21_port, a(20) => PCPlus4F_20_port, 
                           a(19) => PCPlus4F_19_port, a(18) => PCPlus4F_18_port
                           , a(17) => PCPlus4F_17_port, a(16) => 
                           PCPlus4F_16_port, a(15) => PCPlus4F_15_port, a(14) 
                           => PCPlus4F_14_port, a(13) => PCPlus4F_13_port, 
                           a(12) => PCPlus4F_12_port, a(11) => PCPlus4F_11_port
                           , a(10) => PCPlus4F_10_port, a(9) => PCPlus4F_9_port
                           , a(8) => PCPlus4F_8_port, a(7) => PCPlus4F_7_port, 
                           a(6) => PCPlus4F_6_port, a(5) => PCPlus4F_5_port, 
                           a(4) => PCPlus4F_4_port, a(3) => PCPlus4F_3_port, 
                           a(2) => PCPlus4F_2_port, a(1) => PCPlus4F_1_port, 
                           a(0) => PCPlus4F_0_port, b(31) => PCBranchD(31), 
                           b(30) => PCBranchD(30), b(29) => PCBranchD(29), 
                           b(28) => PCBranchD(28), b(27) => PCBranchD(27), 
                           b(26) => PCBranchD(26), b(25) => PCBranchD(25), 
                           b(24) => PCBranchD(24), b(23) => PCBranchD(23), 
                           b(22) => PCBranchD(22), b(21) => PCBranchD(21), 
                           b(20) => PCBranchD(20), b(19) => PCBranchD(19), 
                           b(18) => PCBranchD(18), b(17) => PCBranchD(17), 
                           b(16) => PCBranchD(16), b(15) => PCBranchD(15), 
                           b(14) => PCBranchD(14), b(13) => PCBranchD(13), 
                           b(12) => PCBranchD(12), b(11) => PCBranchD(11), 
                           b(10) => PCBranchD(10), b(9) => PCBranchD(9), b(8) 
                           => PCBranchD(8), b(7) => PCBranchD(7), b(6) => 
                           PCBranchD(6), b(5) => PCBranchD(5), b(4) => 
                           PCBranchD(4), b(3) => PCBranchD(3), b(2) => 
                           PCBranchD(2), b(1) => PCBranchD(1), b(0) => 
                           PCBranchD(0), sel => PCSrcD, y(31) => PC_31_port, 
                           y(30) => PC_30_port, y(29) => PC_29_port, y(28) => 
                           PC_28_port, y(27) => PC_27_port, y(26) => PC_26_port
                           , y(25) => PC_25_port, y(24) => PC_24_port, y(23) =>
                           PC_23_port, y(22) => PC_22_port, y(21) => PC_21_port
                           , y(20) => PC_20_port, y(19) => PC_19_port, y(18) =>
                           PC_18_port, y(17) => PC_17_port, y(16) => PC_16_port
                           , y(15) => PC_15_port, y(14) => PC_14_port, y(13) =>
                           PC_13_port, y(12) => PC_12_port, y(11) => PC_11_port
                           , y(10) => PC_10_port, y(9) => PC_9_port, y(8) => 
                           PC_8_port, y(7) => PC_7_port, y(6) => PC_6_port, 
                           y(5) => PC_5_port, y(4) => PC_4_port, y(3) => 
                           PC_3_port, y(2) => PC_2_port, y(1) => PC_1_port, 
                           y(0) => PC_0_port);
   pc_reg : register_generic_nbit32 port map( d(31) => PC_31_port, d(30) => 
                           PC_30_port, d(29) => PC_29_port, d(28) => PC_28_port
                           , d(27) => PC_27_port, d(26) => PC_26_port, d(25) =>
                           PC_25_port, d(24) => PC_24_port, d(23) => PC_23_port
                           , d(22) => PC_22_port, d(21) => PC_21_port, d(20) =>
                           PC_20_port, d(19) => PC_19_port, d(18) => PC_18_port
                           , d(17) => PC_17_port, d(16) => PC_16_port, d(15) =>
                           PC_15_port, d(14) => PC_14_port, d(13) => PC_13_port
                           , d(12) => PC_12_port, d(11) => PC_11_port, d(10) =>
                           PC_10_port, d(9) => PC_9_port, d(8) => PC_8_port, 
                           d(7) => PC_7_port, d(6) => PC_6_port, d(5) => 
                           PC_5_port, d(4) => PC_4_port, d(3) => PC_3_port, 
                           d(2) => PC_2_port, d(1) => PC_1_port, d(0) => 
                           PC_0_port, q(31) => address_to_iram_31_port, q(30) 
                           => address_to_iram_30_port, q(29) => 
                           address_to_iram_29_port, q(28) => 
                           address_to_iram_28_port, q(27) => 
                           address_to_iram_27_port, q(26) => 
                           address_to_iram_26_port, q(25) => 
                           address_to_iram_25_port, q(24) => 
                           address_to_iram_24_port, q(23) => 
                           address_to_iram_23_port, q(22) => 
                           address_to_iram_22_port, q(21) => 
                           address_to_iram_21_port, q(20) => 
                           address_to_iram_20_port, q(19) => 
                           address_to_iram_19_port, q(18) => 
                           address_to_iram_18_port, q(17) => 
                           address_to_iram_17_port, q(16) => 
                           address_to_iram_16_port, q(15) => 
                           address_to_iram_15_port, q(14) => 
                           address_to_iram_14_port, q(13) => 
                           address_to_iram_13_port, q(12) => 
                           address_to_iram_12_port, q(11) => 
                           address_to_iram_11_port, q(10) => 
                           address_to_iram_10_port, q(9) => 
                           address_to_iram_9_port, q(8) => 
                           address_to_iram_8_port, q(7) => 
                           address_to_iram_7_port, q(6) => 
                           address_to_iram_6_port, q(5) => 
                           address_to_iram_5_port, q(4) => 
                           address_to_iram_4_port, q(3) => 
                           address_to_iram_3_port, q(2) => 
                           address_to_iram_2_port, q(1) => 
                           address_to_iram_1_port, q(0) => 
                           address_to_iram_0_port, clk => clk, reset => rst, en
                           => n1);
   PCPlus4Adder : adder_genericu_nbit32 port map( a(31) => 
                           address_to_iram_31_port, a(30) => 
                           address_to_iram_30_port, a(29) => 
                           address_to_iram_29_port, a(28) => 
                           address_to_iram_28_port, a(27) => 
                           address_to_iram_27_port, a(26) => 
                           address_to_iram_26_port, a(25) => 
                           address_to_iram_25_port, a(24) => 
                           address_to_iram_24_port, a(23) => 
                           address_to_iram_23_port, a(22) => 
                           address_to_iram_22_port, a(21) => 
                           address_to_iram_21_port, a(20) => 
                           address_to_iram_20_port, a(19) => 
                           address_to_iram_19_port, a(18) => 
                           address_to_iram_18_port, a(17) => 
                           address_to_iram_17_port, a(16) => 
                           address_to_iram_16_port, a(15) => 
                           address_to_iram_15_port, a(14) => 
                           address_to_iram_14_port, a(13) => 
                           address_to_iram_13_port, a(12) => 
                           address_to_iram_12_port, a(11) => 
                           address_to_iram_11_port, a(10) => 
                           address_to_iram_10_port, a(9) => 
                           address_to_iram_9_port, a(8) => 
                           address_to_iram_8_port, a(7) => 
                           address_to_iram_7_port, a(6) => 
                           address_to_iram_6_port, a(5) => 
                           address_to_iram_5_port, a(4) => 
                           address_to_iram_4_port, a(3) => 
                           address_to_iram_3_port, a(2) => 
                           address_to_iram_2_port, a(1) => 
                           address_to_iram_1_port, a(0) => 
                           address_to_iram_0_port, b(31) => X_Logic0_port, 
                           b(30) => X_Logic0_port, b(29) => X_Logic0_port, 
                           b(28) => X_Logic0_port, b(27) => X_Logic0_port, 
                           b(26) => X_Logic0_port, b(25) => X_Logic0_port, 
                           b(24) => X_Logic0_port, b(23) => X_Logic0_port, 
                           b(22) => X_Logic0_port, b(21) => X_Logic0_port, 
                           b(20) => X_Logic0_port, b(19) => X_Logic0_port, 
                           b(18) => X_Logic0_port, b(17) => X_Logic0_port, 
                           b(16) => X_Logic0_port, b(15) => X_Logic0_port, 
                           b(14) => X_Logic0_port, b(13) => X_Logic0_port, 
                           b(12) => X_Logic0_port, b(11) => X_Logic0_port, 
                           b(10) => X_Logic0_port, b(9) => X_Logic0_port, b(8) 
                           => X_Logic0_port, b(7) => X_Logic0_port, b(6) => 
                           X_Logic0_port, b(5) => X_Logic0_port, b(4) => 
                           X_Logic0_port, b(3) => X_Logic0_port, b(2) => 
                           X_Logic1_port, b(1) => X_Logic0_port, b(0) => 
                           X_Logic0_port, y(31) => PCPlus4F_31_port, y(30) => 
                           PCPlus4F_30_port, y(29) => PCPlus4F_29_port, y(28) 
                           => PCPlus4F_28_port, y(27) => PCPlus4F_27_port, 
                           y(26) => PCPlus4F_26_port, y(25) => PCPlus4F_25_port
                           , y(24) => PCPlus4F_24_port, y(23) => 
                           PCPlus4F_23_port, y(22) => PCPlus4F_22_port, y(21) 
                           => PCPlus4F_21_port, y(20) => PCPlus4F_20_port, 
                           y(19) => PCPlus4F_19_port, y(18) => PCPlus4F_18_port
                           , y(17) => PCPlus4F_17_port, y(16) => 
                           PCPlus4F_16_port, y(15) => PCPlus4F_15_port, y(14) 
                           => PCPlus4F_14_port, y(13) => PCPlus4F_13_port, 
                           y(12) => PCPlus4F_12_port, y(11) => PCPlus4F_11_port
                           , y(10) => PCPlus4F_10_port, y(9) => PCPlus4F_9_port
                           , y(8) => PCPlus4F_8_port, y(7) => PCPlus4F_7_port, 
                           y(6) => PCPlus4F_6_port, y(5) => PCPlus4F_5_port, 
                           y(4) => PCPlus4F_4_port, y(3) => PCPlus4F_3_port, 
                           y(2) => PCPlus4F_2_port, y(1) => PCPlus4F_1_port, 
                           y(0) => PCPlus4F_0_port);
   U3 : INV_X2 port map( A => StallF, ZN => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity cu is

   port( Rst : in std_logic;  OPCODE : in std_logic_vector (5 downto 0);  FUNC 
         : in std_logic_vector (10 downto 0);  BranchD, Select_ext, IsJal, RD1,
         RD2, RegWriteD : out std_logic;  Comp_control : out std_logic_vector 
         (1 downto 0);  en_ALU, RegDestD, ALUSrcD : out std_logic;  ALUcontrolD
         : out std_logic_vector (5 downto 0);  MemWriteD, MemToRegD, CALL, RET 
         : out std_logic;  FILL, SPILL : in std_logic);

end cu;

architecture SYN_dlx_cu of cu is

signal X_Logic0_port : std_logic;

begin
   BranchD <= X_Logic0_port;
   Select_ext <= X_Logic0_port;
   IsJal <= X_Logic0_port;
   RD1 <= X_Logic0_port;
   RD2 <= X_Logic0_port;
   RegWriteD <= X_Logic0_port;
   Comp_control <= ( X_Logic0_port, X_Logic0_port );
   en_ALU <= X_Logic0_port;
   RegDestD <= X_Logic0_port;
   ALUSrcD <= X_Logic0_port;
   ALUcontrolD <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port,
      X_Logic0_port, X_Logic0_port );
   MemWriteD <= X_Logic0_port;
   MemToRegD <= X_Logic0_port;
   
   X_Logic0_port <= '0';
   RET <= '0';
   CALL <= '0';

end SYN_dlx_cu;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity hazard_detection_unit is

   port( RsD, RtD, RsE, RtE, WriteRegM, WriteRegW, WriteRegE : in 
         std_logic_vector (4 downto 0);  BranchD, MemToRegE, MemToRegM, 
         RegWriteM, RegWriteW, RegWriteE : in std_logic;  ForwardAD, ForwardBD 
         : out std_logic;  ForwardAE, ForwardBE : out std_logic_vector (1 
         downto 0);  StallF, StallD, FlushE : out std_logic);

end hazard_detection_unit;

architecture SYN_behavioral of hazard_detection_unit is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, N15, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13_port, n14, 
      n15_port, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87 : std_logic;

begin
   
   FlushE <= '0';
   U2 : OR3_X1 port map( A1 => n35, A2 => n40, A3 => n41, ZN => N15);
   U3 : INV_X2 port map( A => N15, ZN => ForwardBD);
   U4 : OR3_X1 port map( A1 => n34, A2 => n49, A3 => n41, ZN => N13);
   U5 : INV_X2 port map( A => N13, ZN => ForwardAD);
   U6 : INV_X1 port map( A => n3, ZN => StallF);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => StallD);
   U8 : NAND2_X1 port map( A1 => MemToRegE, A2 => n6, ZN => n3);
   U9 : OAI33_X1 port map( A1 => n7, A2 => n8, A3 => n9, B1 => n10, B2 => n11, 
                           B3 => n12, ZN => n6);
   U10 : XOR2_X1 port map( A => RtE(4), B => RtD(4), Z => n12);
   U11 : XOR2_X1 port map( A => RtE(3), B => RtD(3), Z => n11);
   U12 : NAND3_X1 port map( A1 => n13_port, A2 => n14, A3 => n15_port, ZN => 
                           n10);
   U13 : XNOR2_X1 port map( A => RtD(0), B => RtE(0), ZN => n15_port);
   U14 : XNOR2_X1 port map( A => RtD(1), B => RtE(1), ZN => n14);
   U15 : XNOR2_X1 port map( A => RtD(2), B => RtE(2), ZN => n13_port);
   U16 : XOR2_X1 port map( A => RtE(4), B => RsD(4), Z => n9);
   U17 : XOR2_X1 port map( A => RtE(2), B => RsD(2), Z => n8);
   U18 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => n18, ZN => n7);
   U19 : XNOR2_X1 port map( A => RsD(0), B => RtE(0), ZN => n18);
   U20 : XNOR2_X1 port map( A => RsD(1), B => RtE(1), ZN => n17);
   U21 : XOR2_X1 port map( A => RsD(3), B => n19, Z => n16);
   U22 : INV_X1 port map( A => BranchD, ZN => n5);
   U23 : AOI22_X1 port map( A1 => MemToRegM, A2 => n20, B1 => RegWriteE, B2 => 
                           n21, ZN => n4);
   U24 : OAI33_X1 port map( A1 => n22, A2 => n23, A3 => n24, B1 => n25, B2 => 
                           n26, B3 => n27, ZN => n21);
   U25 : XOR2_X1 port map( A => WriteRegE(4), B => RtD(4), Z => n27);
   U26 : XOR2_X1 port map( A => WriteRegE(3), B => RtD(3), Z => n26);
   U27 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => n25);
   U28 : XNOR2_X1 port map( A => WriteRegE(0), B => RtD(0), ZN => n30);
   U29 : XNOR2_X1 port map( A => WriteRegE(1), B => RtD(1), ZN => n29);
   U30 : XNOR2_X1 port map( A => WriteRegE(2), B => RtD(2), ZN => n28);
   U31 : XOR2_X1 port map( A => WriteRegE(4), B => RsD(4), Z => n24);
   U32 : XOR2_X1 port map( A => WriteRegE(3), B => RsD(3), Z => n23);
   U33 : NAND3_X1 port map( A1 => n31, A2 => n32, A3 => n33, ZN => n22);
   U34 : XNOR2_X1 port map( A => WriteRegE(0), B => RsD(0), ZN => n33);
   U35 : XNOR2_X1 port map( A => WriteRegE(1), B => RsD(1), ZN => n32);
   U36 : XNOR2_X1 port map( A => WriteRegE(2), B => RsD(2), ZN => n31);
   U37 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => n20);
   U38 : NOR2_X1 port map( A1 => n36, A2 => n37, ZN => ForwardBE(1));
   U39 : NOR2_X1 port map( A1 => n38, A2 => n39, ZN => ForwardAE(1));
   U40 : NOR3_X1 port map( A1 => n42, A2 => RtD(1), A3 => RtD(0), ZN => n40);
   U41 : OR3_X1 port map( A1 => RtD(3), A2 => RtD(4), A3 => RtD(2), ZN => n42);
   U42 : NAND4_X1 port map( A1 => n43, A2 => n44, A3 => n45, A4 => n46, ZN => 
                           n35);
   U43 : NOR2_X1 port map( A1 => n47, A2 => n48, ZN => n46);
   U44 : XOR2_X1 port map( A => WriteRegM(4), B => RtD(4), Z => n48);
   U45 : XOR2_X1 port map( A => WriteRegM(3), B => RtD(3), Z => n47);
   U46 : XNOR2_X1 port map( A => RtD(1), B => WriteRegM(1), ZN => n45);
   U47 : XNOR2_X1 port map( A => RtD(2), B => WriteRegM(2), ZN => n44);
   U48 : XNOR2_X1 port map( A => RtD(0), B => WriteRegM(0), ZN => n43);
   U49 : NOR3_X1 port map( A1 => n50, A2 => RsD(1), A3 => RsD(0), ZN => n49);
   U50 : OR3_X1 port map( A1 => RsD(3), A2 => RsD(4), A3 => RsD(2), ZN => n50);
   U51 : NAND4_X1 port map( A1 => n51, A2 => n52, A3 => n53, A4 => n54, ZN => 
                           n34);
   U52 : NOR2_X1 port map( A1 => n55, A2 => n56, ZN => n54);
   U53 : XOR2_X1 port map( A => WriteRegM(4), B => RsD(4), Z => n56);
   U54 : XOR2_X1 port map( A => WriteRegM(3), B => RsD(3), Z => n55);
   U55 : XNOR2_X1 port map( A => RsD(1), B => WriteRegM(1), ZN => n53);
   U56 : XNOR2_X1 port map( A => RsD(2), B => WriteRegM(2), ZN => n52);
   U57 : XNOR2_X1 port map( A => RsD(0), B => WriteRegM(0), ZN => n51);
   U58 : NOR4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           ForwardBE(0));
   U59 : XOR2_X1 port map( A => WriteRegW(3), B => RtE(3), Z => n60);
   U60 : NAND2_X1 port map( A1 => n37, A2 => n61, ZN => n58);
   U61 : INV_X1 port map( A => n36, ZN => n61);
   U62 : NOR4_X1 port map( A1 => RtE(3), A2 => RtE(4), A3 => RtE(2), A4 => n62,
                           ZN => n36);
   U63 : OR2_X1 port map( A1 => RtE(1), A2 => RtE(0), ZN => n62);
   U64 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           n37);
   U65 : NOR3_X1 port map( A1 => n67, A2 => n41, A3 => n68, ZN => n66);
   U66 : XOR2_X1 port map( A => WriteRegM(1), B => RtE(1), Z => n68);
   U67 : XOR2_X1 port map( A => WriteRegM(0), B => RtE(0), Z => n67);
   U68 : XOR2_X1 port map( A => n19, B => WriteRegM(3), Z => n65);
   U69 : INV_X1 port map( A => RtE(3), ZN => n19);
   U70 : XNOR2_X1 port map( A => RtE(4), B => WriteRegM(4), ZN => n64);
   U71 : XNOR2_X1 port map( A => RtE(2), B => WriteRegM(2), ZN => n63);
   U72 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n57);
   U73 : XNOR2_X1 port map( A => WriteRegW(0), B => RtE(0), ZN => n72);
   U74 : XNOR2_X1 port map( A => WriteRegW(1), B => RtE(1), ZN => n71);
   U75 : XNOR2_X1 port map( A => WriteRegW(2), B => RtE(2), ZN => n70);
   U76 : XNOR2_X1 port map( A => WriteRegW(4), B => RtE(4), ZN => n69);
   U77 : NOR4_X1 port map( A1 => n73, A2 => n74, A3 => n59, A4 => n75, ZN => 
                           ForwardAE(0));
   U78 : XOR2_X1 port map( A => WriteRegW(3), B => RsE(3), Z => n75);
   U79 : INV_X1 port map( A => RegWriteW, ZN => n59);
   U80 : NAND2_X1 port map( A1 => n39, A2 => n76, ZN => n74);
   U81 : INV_X1 port map( A => n38, ZN => n76);
   U82 : NOR4_X1 port map( A1 => RsE(3), A2 => RsE(4), A3 => RsE(2), A4 => n77,
                           ZN => n38);
   U83 : OR2_X1 port map( A1 => RsE(1), A2 => RsE(0), ZN => n77);
   U84 : NAND4_X1 port map( A1 => n78, A2 => n79, A3 => n80, A4 => n81, ZN => 
                           n39);
   U85 : NOR3_X1 port map( A1 => n82, A2 => n41, A3 => n83, ZN => n81);
   U86 : XOR2_X1 port map( A => WriteRegM(1), B => RsE(1), Z => n83);
   U87 : INV_X1 port map( A => RegWriteM, ZN => n41);
   U88 : XOR2_X1 port map( A => WriteRegM(0), B => RsE(0), Z => n82);
   U89 : XNOR2_X1 port map( A => RsE(3), B => WriteRegM(3), ZN => n80);
   U90 : XNOR2_X1 port map( A => RsE(4), B => WriteRegM(4), ZN => n79);
   U91 : XNOR2_X1 port map( A => RsE(2), B => WriteRegM(2), ZN => n78);
   U92 : NAND4_X1 port map( A1 => n84, A2 => n85, A3 => n86, A4 => n87, ZN => 
                           n73);
   U93 : XNOR2_X1 port map( A => RsE(0), B => WriteRegW(0), ZN => n87);
   U94 : XNOR2_X1 port map( A => RsE(1), B => WriteRegW(1), ZN => n86);
   U95 : XNOR2_X1 port map( A => RsE(2), B => WriteRegW(2), ZN => n85);
   U96 : XNOR2_X1 port map( A => RsE(4), B => WriteRegW(4), ZN => n84);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity DataPath_wrapper is

   port( clk, rst : in std_logic;  address_to_iram : out std_logic_vector (31 
         downto 0);  iram_to_dlx : in std_logic_vector (31 downto 0);  
         address_to_dram, data_to_dram : out std_logic_vector (31 downto 0);  
         dram_to_dlx : in std_logic_vector (31 downto 0);  dram_we : out 
         std_logic;  StallF, StallD, ForwardAD, ForwardBD, FlushE, rst_RF, 
         en_RF : in std_logic;  RsD_H, RtD_H : out std_logic_vector (4 downto 
         0);  ForwardAE, ForwardBE : in std_logic_vector (1 downto 0);  
         WriteRegE_H, RsE_H, RtE_H, WriteRegMOut_H : out std_logic_vector (4 
         downto 0);  rst_mem : in std_logic;  WriteRegWBOut_H : out 
         std_logic_vector (4 downto 0);  OP : out std_logic_vector (5 downto 0)
         ;  FUNC : out std_logic_vector (10 downto 0);  EqualD, FILL, SPILL : 
         out std_logic;  PCSrcD, RegWriteW, Select_ext, CALL, RET, RD1_EN, 
         RD2_EN, isJal : in std_logic;  Comp_control : in std_logic_vector (1 
         downto 0);  RegDstE, ALUSrcE : in std_logic;  ALUControlE : in 
         std_logic_vector (5 downto 0);  en_ALU, MemWriteM, MemToRegW : in 
         std_logic);

end DataPath_wrapper;

architecture SYN_Behavioral of DataPath_wrapper is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component writeback_unit_N32
      port( ReadDataW, ALUOutW : in std_logic_vector (31 downto 0);  WriteRegW 
            : in std_logic_vector (4 downto 0);  MemToRegW : in std_logic;  
            WriteRegW_out : out std_logic_vector (4 downto 0);  ResultW : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component memory_unit_nbit32_nwords64
      port( ALUOutMIn, WriteDataM : in std_logic_vector (31 downto 0);  
            ReadDataM, ALUOutMOut, address_to_dram, data_to_dram : out 
            std_logic_vector (31 downto 0);  dram_to_dlx : in std_logic_vector 
            (31 downto 0);  WriteRegMIn : in std_logic_vector (4 downto 0);  
            WriteRegMOut : out std_logic_vector (4 downto 0);  clk, rst, 
            MemWriteM : in std_logic;  MemWriteM_out : out std_logic);
   end component;
   
   component execute_stage_wrapper_NBIT32_N32
      port( en_alu : in std_logic;  RD1E, RD2E : in std_logic_vector (31 downto
            0);  RsE, RdE, RtE : in std_logic_vector (4 downto 0);  SignImmE, 
            ALUOutME, ResultWE : in std_logic_vector (31 downto 0);  ALUoutE : 
            out std_logic_vector (31 downto 0);  WriteRegE : out 
            std_logic_vector (4 downto 0);  WriteDataE : out std_logic_vector 
            (31 downto 0);  ForwardAE, ForwardBE : in std_logic_vector (1 
            downto 0);  RsE_o, RtE_o : out std_logic_vector (4 downto 0);  
            RegDstE, ALUSrcE : in std_logic;  ALUcontrolE : in std_logic_vector
            (5 downto 0));
   end component;
   
   component Decode_wrapper
      port( instrD, PcPlus4D : in std_logic_vector (31 downto 0);  select_ext, 
            ForwardAd, ForwardBD, clk, en, rst, RD1_EN, RD2_EN : in std_logic; 
            ALUOutM : in std_logic_vector (31 downto 0);  WriteRegW : in 
            std_logic_vector (4 downto 0);  ResultW : in std_logic_vector (31 
            downto 0);  CALL, RET, IsJal : in std_logic;  Comp_control : in 
            std_logic_vector (1 downto 0);  RegWriteW : in std_logic;  
            Memory_in : in std_logic_vector (31 downto 0);  Memory_out : out 
            std_logic_vector (31 downto 0);  FILL, SPILL : out std_logic;  RsD,
            RtD, RdE : out std_logic_vector (4 downto 0);  SignImmD, PCBranchD 
            : out std_logic_vector (31 downto 0);  EqualD : out std_logic;  OP 
            : out std_logic_vector (5 downto 0);  FUNC : out std_logic_vector 
            (10 downto 0);  RD1, RD2 : out std_logic_vector (31 downto 0));
   end component;
   
   component fetch_stage_wrapper_nbit32_nwords64
      port( PCBranchD : in std_logic_vector (31 downto 0);  PCPlus4F, InstrD, 
            address_to_iram : out std_logic_vector (31 downto 0);  iram_to_dlx 
            : in std_logic_vector (31 downto 0);  PCSrcD, StallF, clk, rst : in
            std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, RsD_H_4_port, RsD_H_3_port, RsD_H_2_port, RsD_H_1_port
      , RsD_H_0_port, RtD_H_4_port, RtD_H_3_port, RtD_H_2_port, RtD_H_1_port, 
      RtD_H_0_port, WriteRegE_H_4_port, WriteRegE_H_3_port, WriteRegE_H_2_port,
      WriteRegE_H_1_port, WriteRegE_H_0_port, WriteRegMOut_H_4_port, 
      WriteRegMOut_H_3_port, WriteRegMOut_H_2_port, WriteRegMOut_H_1_port, 
      WriteRegMOut_H_0_port, WriteRegWBOut_H_4_port, WriteRegWBOut_H_3_port, 
      WriteRegWBOut_H_2_port, WriteRegWBOut_H_1_port, WriteRegWBOut_H_0_port, 
      IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, IR_26_port, 
      IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, IR_20_port, 
      IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, IR_14_port, 
      IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, IR_8_port, 
      IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, IR_2_port, 
      IR_1_port, IR_0_port, PCPlus4_31_port, PCPlus4_30_port, PCPlus4_29_port, 
      PCPlus4_28_port, PCPlus4_27_port, PCPlus4_26_port, PCPlus4_25_port, 
      PCPlus4_24_port, PCPlus4_23_port, PCPlus4_22_port, PCPlus4_21_port, 
      PCPlus4_20_port, PCPlus4_19_port, PCPlus4_18_port, PCPlus4_17_port, 
      PCPlus4_16_port, PCPlus4_15_port, PCPlus4_14_port, PCPlus4_13_port, 
      PCPlus4_12_port, PCPlus4_11_port, PCPlus4_10_port, PCPlus4_9_port, 
      PCPlus4_8_port, PCPlus4_7_port, PCPlus4_6_port, PCPlus4_5_port, 
      PCPlus4_4_port, PCPlus4_3_port, PCPlus4_2_port, PCPlus4_1_port, 
      PCPlus4_0_port, RD1_31_port, RD1_30_port, RD1_29_port, RD1_28_port, 
      RD1_27_port, RD1_26_port, RD1_25_port, RD1_24_port, RD1_23_port, 
      RD1_22_port, RD1_21_port, RD1_20_port, RD1_19_port, RD1_18_port, 
      RD1_17_port, RD1_16_port, RD1_15_port, RD1_14_port, RD1_13_port, 
      RD1_12_port, RD1_11_port, RD1_10_port, RD1_9_port, RD1_8_port, RD1_7_port
      , RD1_6_port, RD1_5_port, RD1_4_port, RD1_3_port, RD1_2_port, RD1_1_port,
      RD1_0_port, RD2_31_port, RD2_30_port, RD2_29_port, RD2_28_port, 
      RD2_27_port, RD2_26_port, RD2_25_port, RD2_24_port, RD2_23_port, 
      RD2_22_port, RD2_21_port, RD2_20_port, RD2_19_port, RD2_18_port, 
      RD2_17_port, RD2_16_port, RD2_15_port, RD2_14_port, RD2_13_port, 
      RD2_12_port, RD2_11_port, RD2_10_port, RD2_9_port, RD2_8_port, RD2_7_port
      , RD2_6_port, RD2_5_port, RD2_4_port, RD2_3_port, RD2_2_port, RD2_1_port,
      RD2_0_port, RsD_4_port, RsD_3_port, RsD_2_port, RsD_1_port, RsD_0_port, 
      RtD_4_port, RtD_3_port, RtD_2_port, RtD_1_port, RtD_0_port, RdD_4_port, 
      RdD_3_port, RdD_2_port, RdD_1_port, RdD_0_port, SignImmD_31_port, 
      SignImmD_30_port, SignImmD_29_port, SignImmD_28_port, SignImmD_27_port, 
      SignImmD_26_port, SignImmD_25_port, SignImmD_24_port, SignImmD_23_port, 
      SignImmD_22_port, SignImmD_21_port, SignImmD_20_port, SignImmD_19_port, 
      SignImmD_18_port, SignImmD_17_port, SignImmD_16_port, SignImmD_15_port, 
      SignImmD_14_port, SignImmD_13_port, SignImmD_12_port, SignImmD_11_port, 
      SignImmD_10_port, SignImmD_9_port, SignImmD_8_port, SignImmD_7_port, 
      SignImmD_6_port, SignImmD_5_port, SignImmD_4_port, SignImmD_3_port, 
      SignImmD_2_port, SignImmD_1_port, SignImmD_0_port, ALUOutE_31_port, 
      ALUOutE_30_port, ALUOutE_29_port, ALUOutE_28_port, ALUOutE_27_port, 
      ALUOutE_26_port, ALUOutE_25_port, ALUOutE_24_port, ALUOutE_23_port, 
      ALUOutE_22_port, ALUOutE_21_port, ALUOutE_20_port, ALUOutE_19_port, 
      ALUOutE_18_port, ALUOutE_17_port, ALUOutE_16_port, ALUOutE_15_port, 
      ALUOutE_14_port, ALUOutE_13_port, ALUOutE_12_port, ALUOutE_11_port, 
      ALUOutE_10_port, ALUOutE_9_port, ALUOutE_8_port, ALUOutE_7_port, 
      ALUOutE_6_port, ALUOutE_5_port, ALUOutE_4_port, ALUOutE_3_port, 
      ALUOutE_2_port, ALUOutE_1_port, ALUOutE_0_port, WriteDataE_31_port, 
      WriteDataE_30_port, WriteDataE_29_port, WriteDataE_28_port, 
      WriteDataE_27_port, WriteDataE_26_port, WriteDataE_25_port, 
      WriteDataE_24_port, WriteDataE_23_port, WriteDataE_22_port, 
      WriteDataE_21_port, WriteDataE_20_port, WriteDataE_19_port, 
      WriteDataE_18_port, WriteDataE_17_port, WriteDataE_16_port, 
      WriteDataE_15_port, WriteDataE_14_port, WriteDataE_13_port, 
      WriteDataE_12_port, WriteDataE_11_port, WriteDataE_10_port, 
      WriteDataE_9_port, WriteDataE_8_port, WriteDataE_7_port, 
      WriteDataE_6_port, WriteDataE_5_port, WriteDataE_4_port, 
      WriteDataE_3_port, WriteDataE_2_port, WriteDataE_1_port, 
      WriteDataE_0_port, WriteRegE_4_port, WriteRegE_3_port, WriteRegE_2_port, 
      WriteRegE_1_port, WriteRegE_0_port, ReadDataM_31_port, ReadDataM_30_port,
      ReadDataM_29_port, ReadDataM_28_port, ReadDataM_27_port, 
      ReadDataM_26_port, ReadDataM_25_port, ReadDataM_24_port, 
      ReadDataM_23_port, ReadDataM_22_port, ReadDataM_21_port, 
      ReadDataM_20_port, ReadDataM_19_port, ReadDataM_18_port, 
      ReadDataM_17_port, ReadDataM_16_port, ReadDataM_15_port, 
      ReadDataM_14_port, ReadDataM_13_port, ReadDataM_12_port, 
      ReadDataM_11_port, ReadDataM_10_port, ReadDataM_9_port, ReadDataM_8_port,
      ReadDataM_7_port, ReadDataM_6_port, ReadDataM_5_port, ReadDataM_4_port, 
      ReadDataM_3_port, ReadDataM_2_port, ReadDataM_1_port, ReadDataM_0_port, 
      ALUOutM_31_port, ALUOutM_30_port, ALUOutM_29_port, ALUOutM_28_port, 
      ALUOutM_27_port, ALUOutM_26_port, ALUOutM_25_port, ALUOutM_24_port, 
      ALUOutM_23_port, ALUOutM_22_port, ALUOutM_21_port, ALUOutM_20_port, 
      ALUOutM_19_port, ALUOutM_18_port, ALUOutM_17_port, ALUOutM_16_port, 
      ALUOutM_15_port, ALUOutM_14_port, ALUOutM_13_port, ALUOutM_12_port, 
      ALUOutM_11_port, ALUOutM_10_port, ALUOutM_9_port, ALUOutM_8_port, 
      ALUOutM_7_port, ALUOutM_6_port, ALUOutM_5_port, ALUOutM_4_port, 
      ALUOutM_3_port, ALUOutM_2_port, ALUOutM_1_port, ALUOutM_0_port, 
      WriteRegM_4_port, WriteRegM_3_port, WriteRegM_2_port, WriteRegM_1_port, 
      WriteRegM_0_port, PCBranchD_wire_31_port, PCBranchD_wire_30_port, 
      PCBranchD_wire_29_port, PCBranchD_wire_28_port, PCBranchD_wire_27_port, 
      PCBranchD_wire_26_port, PCBranchD_wire_25_port, PCBranchD_wire_24_port, 
      PCBranchD_wire_23_port, PCBranchD_wire_22_port, PCBranchD_wire_21_port, 
      PCBranchD_wire_20_port, PCBranchD_wire_19_port, PCBranchD_wire_18_port, 
      PCBranchD_wire_17_port, PCBranchD_wire_16_port, PCBranchD_wire_15_port, 
      PCBranchD_wire_14_port, PCBranchD_wire_13_port, PCBranchD_wire_12_port, 
      PCBranchD_wire_11_port, PCBranchD_wire_10_port, PCBranchD_wire_9_port, 
      PCBranchD_wire_8_port, PCBranchD_wire_7_port, PCBranchD_wire_6_port, 
      PCBranchD_wire_5_port, PCBranchD_wire_4_port, PCBranchD_wire_3_port, 
      PCBranchD_wire_2_port, PCBranchD_wire_1_port, PCBranchD_wire_0_port, 
      PCPlus4F_wire_31_port, PCPlus4F_wire_30_port, PCPlus4F_wire_29_port, 
      PCPlus4F_wire_28_port, PCPlus4F_wire_27_port, PCPlus4F_wire_26_port, 
      PCPlus4F_wire_25_port, PCPlus4F_wire_24_port, PCPlus4F_wire_23_port, 
      PCPlus4F_wire_22_port, PCPlus4F_wire_21_port, PCPlus4F_wire_20_port, 
      PCPlus4F_wire_19_port, PCPlus4F_wire_18_port, PCPlus4F_wire_17_port, 
      PCPlus4F_wire_16_port, PCPlus4F_wire_15_port, PCPlus4F_wire_14_port, 
      PCPlus4F_wire_13_port, PCPlus4F_wire_12_port, PCPlus4F_wire_11_port, 
      PCPlus4F_wire_10_port, PCPlus4F_wire_9_port, PCPlus4F_wire_8_port, 
      PCPlus4F_wire_7_port, PCPlus4F_wire_6_port, PCPlus4F_wire_5_port, 
      PCPlus4F_wire_4_port, PCPlus4F_wire_3_port, PCPlus4F_wire_2_port, 
      PCPlus4F_wire_1_port, PCPlus4F_wire_0_port, InstrD_wire_31_port, 
      InstrD_wire_30_port, InstrD_wire_29_port, InstrD_wire_28_port, 
      InstrD_wire_27_port, InstrD_wire_26_port, InstrD_wire_25_port, 
      InstrD_wire_24_port, InstrD_wire_23_port, InstrD_wire_22_port, 
      InstrD_wire_21_port, InstrD_wire_20_port, InstrD_wire_19_port, 
      InstrD_wire_18_port, InstrD_wire_17_port, InstrD_wire_16_port, 
      InstrD_wire_15_port, InstrD_wire_14_port, InstrD_wire_13_port, 
      InstrD_wire_12_port, InstrD_wire_11_port, InstrD_wire_10_port, 
      InstrD_wire_9_port, InstrD_wire_8_port, InstrD_wire_7_port, 
      InstrD_wire_6_port, InstrD_wire_5_port, InstrD_wire_4_port, 
      InstrD_wire_3_port, InstrD_wire_2_port, InstrD_wire_1_port, 
      InstrD_wire_0_port, ALUOutMOut_wire_31_port, ALUOutMOut_wire_30_port, 
      ALUOutMOut_wire_29_port, ALUOutMOut_wire_28_port, ALUOutMOut_wire_27_port
      , ALUOutMOut_wire_26_port, ALUOutMOut_wire_25_port, 
      ALUOutMOut_wire_24_port, ALUOutMOut_wire_23_port, ALUOutMOut_wire_22_port
      , ALUOutMOut_wire_21_port, ALUOutMOut_wire_20_port, 
      ALUOutMOut_wire_19_port, ALUOutMOut_wire_18_port, ALUOutMOut_wire_17_port
      , ALUOutMOut_wire_16_port, ALUOutMOut_wire_15_port, 
      ALUOutMOut_wire_14_port, ALUOutMOut_wire_13_port, ALUOutMOut_wire_12_port
      , ALUOutMOut_wire_11_port, ALUOutMOut_wire_10_port, 
      ALUOutMOut_wire_9_port, ALUOutMOut_wire_8_port, ALUOutMOut_wire_7_port, 
      ALUOutMOut_wire_6_port, ALUOutMOut_wire_5_port, ALUOutMOut_wire_4_port, 
      ALUOutMOut_wire_3_port, ALUOutMOut_wire_2_port, ALUOutMOut_wire_1_port, 
      ALUOutMOut_wire_0_port, ResultW_wire_31_port, ResultW_wire_30_port, 
      ResultW_wire_29_port, ResultW_wire_28_port, ResultW_wire_27_port, 
      ResultW_wire_26_port, ResultW_wire_25_port, ResultW_wire_24_port, 
      ResultW_wire_23_port, ResultW_wire_22_port, ResultW_wire_21_port, 
      ResultW_wire_20_port, ResultW_wire_19_port, ResultW_wire_18_port, 
      ResultW_wire_17_port, ResultW_wire_16_port, ResultW_wire_15_port, 
      ResultW_wire_14_port, ResultW_wire_13_port, ResultW_wire_12_port, 
      ResultW_wire_11_port, ResultW_wire_10_port, ResultW_wire_9_port, 
      ResultW_wire_8_port, ResultW_wire_7_port, ResultW_wire_6_port, 
      ResultW_wire_5_port, ResultW_wire_4_port, ResultW_wire_3_port, 
      ResultW_wire_2_port, ResultW_wire_1_port, ResultW_wire_0_port, 
      RdD_wire_4_port, RdD_wire_3_port, RdD_wire_2_port, RdD_wire_1_port, 
      RdD_wire_0_port, SignImmD_wire_31_port, SignImmD_wire_30_port, 
      SignImmD_wire_29_port, SignImmD_wire_28_port, SignImmD_wire_27_port, 
      SignImmD_wire_26_port, SignImmD_wire_25_port, SignImmD_wire_24_port, 
      SignImmD_wire_23_port, SignImmD_wire_22_port, SignImmD_wire_21_port, 
      SignImmD_wire_20_port, SignImmD_wire_19_port, SignImmD_wire_18_port, 
      SignImmD_wire_17_port, SignImmD_wire_16_port, SignImmD_wire_15_port, 
      SignImmD_wire_14_port, SignImmD_wire_13_port, SignImmD_wire_12_port, 
      SignImmD_wire_11_port, SignImmD_wire_10_port, SignImmD_wire_9_port, 
      SignImmD_wire_8_port, SignImmD_wire_7_port, SignImmD_wire_6_port, 
      SignImmD_wire_5_port, SignImmD_wire_4_port, SignImmD_wire_3_port, 
      SignImmD_wire_2_port, SignImmD_wire_1_port, SignImmD_wire_0_port, 
      RD1_wire_31_port, RD1_wire_30_port, RD1_wire_29_port, RD1_wire_28_port, 
      RD1_wire_27_port, RD1_wire_26_port, RD1_wire_25_port, RD1_wire_24_port, 
      RD1_wire_23_port, RD1_wire_22_port, RD1_wire_21_port, RD1_wire_20_port, 
      RD1_wire_19_port, RD1_wire_18_port, RD1_wire_17_port, RD1_wire_16_port, 
      RD1_wire_15_port, RD1_wire_14_port, RD1_wire_13_port, RD1_wire_12_port, 
      RD1_wire_11_port, RD1_wire_10_port, RD1_wire_9_port, RD1_wire_8_port, 
      RD1_wire_7_port, RD1_wire_6_port, RD1_wire_5_port, RD1_wire_4_port, 
      RD1_wire_3_port, RD1_wire_2_port, RD1_wire_1_port, RD1_wire_0_port, 
      RD2_wire_31_port, RD2_wire_30_port, RD2_wire_29_port, RD2_wire_28_port, 
      RD2_wire_27_port, RD2_wire_26_port, RD2_wire_25_port, RD2_wire_24_port, 
      RD2_wire_23_port, RD2_wire_22_port, RD2_wire_21_port, RD2_wire_20_port, 
      RD2_wire_19_port, RD2_wire_18_port, RD2_wire_17_port, RD2_wire_16_port, 
      RD2_wire_15_port, RD2_wire_14_port, RD2_wire_13_port, RD2_wire_12_port, 
      RD2_wire_11_port, RD2_wire_10_port, RD2_wire_9_port, RD2_wire_8_port, 
      RD2_wire_7_port, RD2_wire_6_port, RD2_wire_5_port, RD2_wire_4_port, 
      RD2_wire_3_port, RD2_wire_2_port, RD2_wire_1_port, RD2_wire_0_port, 
      ALUOutE_wire_31_port, ALUOutE_wire_30_port, ALUOutE_wire_29_port, 
      ALUOutE_wire_28_port, ALUOutE_wire_27_port, ALUOutE_wire_26_port, 
      ALUOutE_wire_25_port, ALUOutE_wire_24_port, ALUOutE_wire_23_port, 
      ALUOutE_wire_22_port, ALUOutE_wire_21_port, ALUOutE_wire_20_port, 
      ALUOutE_wire_19_port, ALUOutE_wire_18_port, ALUOutE_wire_17_port, 
      ALUOutE_wire_16_port, ALUOutE_wire_15_port, ALUOutE_wire_14_port, 
      ALUOutE_wire_13_port, ALUOutE_wire_12_port, ALUOutE_wire_11_port, 
      ALUOutE_wire_10_port, ALUOutE_wire_9_port, ALUOutE_wire_8_port, 
      ALUOutE_wire_7_port, ALUOutE_wire_6_port, ALUOutE_wire_5_port, 
      ALUOutE_wire_4_port, ALUOutE_wire_3_port, ALUOutE_wire_2_port, 
      ALUOutE_wire_1_port, ALUOutE_wire_0_port, WriteDataE_wire_31_port, 
      WriteDataE_wire_30_port, WriteDataE_wire_29_port, WriteDataE_wire_28_port
      , WriteDataE_wire_27_port, WriteDataE_wire_26_port, 
      WriteDataE_wire_25_port, WriteDataE_wire_24_port, WriteDataE_wire_23_port
      , WriteDataE_wire_22_port, WriteDataE_wire_21_port, 
      WriteDataE_wire_20_port, WriteDataE_wire_19_port, WriteDataE_wire_18_port
      , WriteDataE_wire_17_port, WriteDataE_wire_16_port, 
      WriteDataE_wire_15_port, WriteDataE_wire_14_port, WriteDataE_wire_13_port
      , WriteDataE_wire_12_port, WriteDataE_wire_11_port, 
      WriteDataE_wire_10_port, WriteDataE_wire_9_port, WriteDataE_wire_8_port, 
      WriteDataE_wire_7_port, WriteDataE_wire_6_port, WriteDataE_wire_5_port, 
      WriteDataE_wire_4_port, WriteDataE_wire_3_port, WriteDataE_wire_2_port, 
      WriteDataE_wire_1_port, WriteDataE_wire_0_port, ReadDataM_wire_31_port, 
      ReadDataM_wire_30_port, ReadDataM_wire_29_port, ReadDataM_wire_28_port, 
      ReadDataM_wire_27_port, ReadDataM_wire_26_port, ReadDataM_wire_25_port, 
      ReadDataM_wire_24_port, ReadDataM_wire_23_port, ReadDataM_wire_22_port, 
      ReadDataM_wire_21_port, ReadDataM_wire_20_port, ReadDataM_wire_19_port, 
      ReadDataM_wire_18_port, ReadDataM_wire_17_port, ReadDataM_wire_16_port, 
      ReadDataM_wire_15_port, ReadDataM_wire_14_port, ReadDataM_wire_13_port, 
      ReadDataM_wire_12_port, ReadDataM_wire_11_port, ReadDataM_wire_10_port, 
      ReadDataM_wire_9_port, ReadDataM_wire_8_port, ReadDataM_wire_7_port, 
      ReadDataM_wire_6_port, ReadDataM_wire_5_port, ReadDataM_wire_4_port, 
      ReadDataM_wire_3_port, ReadDataM_wire_2_port, ReadDataM_wire_1_port, 
      ReadDataM_wire_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, 
      n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, 
      n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, 
      n_1826, n_1827, n_1828, n_1829, n_1830 : std_logic;

begin
   RsD_H <= ( RsD_H_4_port, RsD_H_3_port, RsD_H_2_port, RsD_H_1_port, 
      RsD_H_0_port );
   RtD_H <= ( RtD_H_4_port, RtD_H_3_port, RtD_H_2_port, RtD_H_1_port, 
      RtD_H_0_port );
   WriteRegE_H <= ( WriteRegE_H_4_port, WriteRegE_H_3_port, WriteRegE_H_2_port,
      WriteRegE_H_1_port, WriteRegE_H_0_port );
   WriteRegMOut_H <= ( WriteRegMOut_H_4_port, WriteRegMOut_H_3_port, 
      WriteRegMOut_H_2_port, WriteRegMOut_H_1_port, WriteRegMOut_H_0_port );
   WriteRegWBOut_H <= ( WriteRegWBOut_H_4_port, WriteRegWBOut_H_3_port, 
      WriteRegWBOut_H_2_port, WriteRegWBOut_H_1_port, WriteRegWBOut_H_0_port );
   
   X_Logic0_port <= '0';
   ALUOutM_reg_0_inst : DFFR_X1 port map( D => ALUOutMOut_wire_0_port, CK => 
                           clk, RN => n14, Q => ALUOutM_0_port, QN => n_1549);
   RD2_reg_0_inst : DFFR_X1 port map( D => RD2_wire_0_port, CK => clk, RN => 
                           n14, Q => RD2_0_port, QN => n_1550);
   RD2_reg_1_inst : DFFR_X1 port map( D => RD2_wire_1_port, CK => clk, RN => n1
                           , Q => RD2_1_port, QN => n_1551);
   RD2_reg_2_inst : DFFR_X1 port map( D => RD2_wire_2_port, CK => clk, RN => n1
                           , Q => RD2_2_port, QN => n_1552);
   RD2_reg_3_inst : DFFR_X1 port map( D => RD2_wire_3_port, CK => clk, RN => n2
                           , Q => RD2_3_port, QN => n_1553);
   RD2_reg_4_inst : DFFR_X1 port map( D => RD2_wire_4_port, CK => clk, RN => 
                           n13, Q => RD2_4_port, QN => n_1554);
   RD2_reg_5_inst : DFFR_X1 port map( D => RD2_wire_5_port, CK => clk, RN => n5
                           , Q => RD2_5_port, QN => n_1555);
   RD2_reg_6_inst : DFFR_X1 port map( D => RD2_wire_6_port, CK => clk, RN => n2
                           , Q => RD2_6_port, QN => n_1556);
   RD2_reg_7_inst : DFFR_X1 port map( D => RD2_wire_7_port, CK => clk, RN => n2
                           , Q => RD2_7_port, QN => n_1557);
   RD2_reg_8_inst : DFFR_X1 port map( D => RD2_wire_8_port, CK => clk, RN => n5
                           , Q => RD2_8_port, QN => n_1558);
   RD2_reg_9_inst : DFFR_X1 port map( D => RD2_wire_9_port, CK => clk, RN => 
                           n12, Q => RD2_9_port, QN => n_1559);
   RD2_reg_10_inst : DFFR_X1 port map( D => RD2_wire_10_port, CK => clk, RN => 
                           n3, Q => RD2_10_port, QN => n_1560);
   RD2_reg_11_inst : DFFR_X1 port map( D => RD2_wire_11_port, CK => clk, RN => 
                           n4, Q => RD2_11_port, QN => n_1561);
   RD2_reg_12_inst : DFFR_X1 port map( D => RD2_wire_12_port, CK => clk, RN => 
                           n11, Q => RD2_12_port, QN => n_1562);
   RD2_reg_13_inst : DFFR_X1 port map( D => RD2_wire_13_port, CK => clk, RN => 
                           n3, Q => RD2_13_port, QN => n_1563);
   RD2_reg_14_inst : DFFR_X1 port map( D => RD2_wire_14_port, CK => clk, RN => 
                           n4, Q => RD2_14_port, QN => n_1564);
   RD2_reg_15_inst : DFFR_X1 port map( D => RD2_wire_15_port, CK => clk, RN => 
                           n6, Q => RD2_15_port, QN => n_1565);
   RD2_reg_16_inst : DFFR_X1 port map( D => RD2_wire_16_port, CK => clk, RN => 
                           n13, Q => RD2_16_port, QN => n_1566);
   RD2_reg_17_inst : DFFR_X1 port map( D => RD2_wire_17_port, CK => clk, RN => 
                           n7, Q => RD2_17_port, QN => n_1567);
   RD2_reg_18_inst : DFFR_X1 port map( D => RD2_wire_18_port, CK => clk, RN => 
                           n7, Q => RD2_18_port, QN => n_1568);
   RD2_reg_19_inst : DFFR_X1 port map( D => RD2_wire_19_port, CK => clk, RN => 
                           n7, Q => RD2_19_port, QN => n_1569);
   RD2_reg_20_inst : DFFR_X1 port map( D => RD2_wire_20_port, CK => clk, RN => 
                           n8, Q => RD2_20_port, QN => n_1570);
   RD2_reg_21_inst : DFFR_X1 port map( D => RD2_wire_21_port, CK => clk, RN => 
                           n8, Q => RD2_21_port, QN => n_1571);
   RD2_reg_22_inst : DFFR_X1 port map( D => RD2_wire_22_port, CK => clk, RN => 
                           n9, Q => RD2_22_port, QN => n_1572);
   RD2_reg_23_inst : DFFR_X1 port map( D => RD2_wire_23_port, CK => clk, RN => 
                           n9, Q => RD2_23_port, QN => n_1573);
   RD2_reg_24_inst : DFFR_X1 port map( D => RD2_wire_24_port, CK => clk, RN => 
                           n11, Q => RD2_24_port, QN => n_1574);
   RD2_reg_25_inst : DFFR_X1 port map( D => RD2_wire_25_port, CK => clk, RN => 
                           n10, Q => RD2_25_port, QN => n_1575);
   RD2_reg_26_inst : DFFR_X1 port map( D => RD2_wire_26_port, CK => clk, RN => 
                           n10, Q => RD2_26_port, QN => n_1576);
   RD2_reg_27_inst : DFFR_X1 port map( D => RD2_wire_27_port, CK => clk, RN => 
                           n10, Q => RD2_27_port, QN => n_1577);
   RD2_reg_28_inst : DFFR_X1 port map( D => RD2_wire_28_port, CK => clk, RN => 
                           n12, Q => RD2_28_port, QN => n_1578);
   RD2_reg_29_inst : DFFR_X1 port map( D => RD2_wire_29_port, CK => clk, RN => 
                           n5, Q => RD2_29_port, QN => n_1579);
   RD2_reg_30_inst : DFFR_X1 port map( D => RD2_wire_30_port, CK => clk, RN => 
                           n6, Q => RD2_30_port, QN => n_1580);
   RD2_reg_31_inst : DFFR_X1 port map( D => RD2_wire_31_port, CK => clk, RN => 
                           n12, Q => RD2_31_port, QN => n_1581);
   RD1_reg_0_inst : DFFR_X1 port map( D => RD1_wire_0_port, CK => clk, RN => 
                           n14, Q => RD1_0_port, QN => n_1582);
   RD1_reg_1_inst : DFFR_X1 port map( D => RD1_wire_1_port, CK => clk, RN => n1
                           , Q => RD1_1_port, QN => n_1583);
   RD1_reg_2_inst : DFFR_X1 port map( D => RD1_wire_2_port, CK => clk, RN => n1
                           , Q => RD1_2_port, QN => n_1584);
   RD1_reg_3_inst : DFFR_X1 port map( D => RD1_wire_3_port, CK => clk, RN => n1
                           , Q => RD1_3_port, QN => n_1585);
   RD1_reg_4_inst : DFFR_X1 port map( D => RD1_wire_4_port, CK => clk, RN => 
                           n13, Q => RD1_4_port, QN => n_1586);
   RD1_reg_5_inst : DFFR_X1 port map( D => RD1_wire_5_port, CK => clk, RN => n5
                           , Q => RD1_5_port, QN => n_1587);
   RD1_reg_6_inst : DFFR_X1 port map( D => RD1_wire_6_port, CK => clk, RN => n2
                           , Q => RD1_6_port, QN => n_1588);
   RD1_reg_7_inst : DFFR_X1 port map( D => RD1_wire_7_port, CK => clk, RN => n2
                           , Q => RD1_7_port, QN => n_1589);
   RD1_reg_8_inst : DFFR_X1 port map( D => RD1_wire_8_port, CK => clk, RN => n4
                           , Q => RD1_8_port, QN => n_1590);
   RD1_reg_9_inst : DFFR_X1 port map( D => RD1_wire_9_port, CK => clk, RN => 
                           n11, Q => RD1_9_port, QN => n_1591);
   RD1_reg_10_inst : DFFR_X1 port map( D => RD1_wire_10_port, CK => clk, RN => 
                           n3, Q => RD1_10_port, QN => n_1592);
   RD1_reg_11_inst : DFFR_X1 port map( D => RD1_wire_11_port, CK => clk, RN => 
                           n4, Q => RD1_11_port, QN => n_1593);
   RD1_reg_12_inst : DFFR_X1 port map( D => RD1_wire_12_port, CK => clk, RN => 
                           n11, Q => RD1_12_port, QN => n_1594);
   RD1_reg_13_inst : DFFR_X1 port map( D => RD1_wire_13_port, CK => clk, RN => 
                           n3, Q => RD1_13_port, QN => n_1595);
   RD1_reg_14_inst : DFFR_X1 port map( D => RD1_wire_14_port, CK => clk, RN => 
                           n4, Q => RD1_14_port, QN => n_1596);
   RD1_reg_15_inst : DFFR_X1 port map( D => RD1_wire_15_port, CK => clk, RN => 
                           n6, Q => RD1_15_port, QN => n_1597);
   RD1_reg_16_inst : DFFR_X1 port map( D => RD1_wire_16_port, CK => clk, RN => 
                           n13, Q => RD1_16_port, QN => n_1598);
   RD1_reg_17_inst : DFFR_X1 port map( D => RD1_wire_17_port, CK => clk, RN => 
                           n6, Q => RD1_17_port, QN => n_1599);
   RD1_reg_18_inst : DFFR_X1 port map( D => RD1_wire_18_port, CK => clk, RN => 
                           n7, Q => RD1_18_port, QN => n_1600);
   RD1_reg_19_inst : DFFR_X1 port map( D => RD1_wire_19_port, CK => clk, RN => 
                           n7, Q => RD1_19_port, QN => n_1601);
   RD1_reg_20_inst : DFFR_X1 port map( D => RD1_wire_20_port, CK => clk, RN => 
                           n8, Q => RD1_20_port, QN => n_1602);
   RD1_reg_21_inst : DFFR_X1 port map( D => RD1_wire_21_port, CK => clk, RN => 
                           n8, Q => RD1_21_port, QN => n_1603);
   RD1_reg_22_inst : DFFR_X1 port map( D => RD1_wire_22_port, CK => clk, RN => 
                           n9, Q => RD1_22_port, QN => n_1604);
   RD1_reg_23_inst : DFFR_X1 port map( D => RD1_wire_23_port, CK => clk, RN => 
                           n9, Q => RD1_23_port, QN => n_1605);
   RD1_reg_24_inst : DFFR_X1 port map( D => RD1_wire_24_port, CK => clk, RN => 
                           n11, Q => RD1_24_port, QN => n_1606);
   RD1_reg_25_inst : DFFR_X1 port map( D => RD1_wire_25_port, CK => clk, RN => 
                           n9, Q => RD1_25_port, QN => n_1607);
   RD1_reg_26_inst : DFFR_X1 port map( D => RD1_wire_26_port, CK => clk, RN => 
                           n10, Q => RD1_26_port, QN => n_1608);
   RD1_reg_27_inst : DFFR_X1 port map( D => RD1_wire_27_port, CK => clk, RN => 
                           n10, Q => RD1_27_port, QN => n_1609);
   RD1_reg_28_inst : DFFR_X1 port map( D => RD1_wire_28_port, CK => clk, RN => 
                           n12, Q => RD1_28_port, QN => n_1610);
   RD1_reg_29_inst : DFFR_X1 port map( D => RD1_wire_29_port, CK => clk, RN => 
                           n5, Q => RD1_29_port, QN => n_1611);
   RD1_reg_30_inst : DFFR_X1 port map( D => RD1_wire_30_port, CK => clk, RN => 
                           n6, Q => RD1_30_port, QN => n_1612);
   RD1_reg_31_inst : DFFR_X1 port map( D => RD1_wire_31_port, CK => clk, RN => 
                           n12, Q => RD1_31_port, QN => n_1613);
   IR_reg_0_inst : DFFR_X1 port map( D => n190, CK => clk, RN => n17, Q => 
                           IR_0_port, QN => n157);
   IR_reg_1_inst : DFFR_X1 port map( D => n191, CK => clk, RN => n17, Q => 
                           IR_1_port, QN => n156);
   IR_reg_2_inst : DFFR_X1 port map( D => n192, CK => clk, RN => n17, Q => 
                           IR_2_port, QN => n155);
   IR_reg_3_inst : DFFR_X1 port map( D => n193, CK => clk, RN => n17, Q => 
                           IR_3_port, QN => n154);
   IR_reg_4_inst : DFFR_X1 port map( D => n194, CK => clk, RN => n17, Q => 
                           IR_4_port, QN => n153);
   IR_reg_5_inst : DFFR_X1 port map( D => n195, CK => clk, RN => n17, Q => 
                           IR_5_port, QN => n152);
   IR_reg_6_inst : DFFR_X1 port map( D => n196, CK => clk, RN => n18, Q => 
                           IR_6_port, QN => n151);
   IR_reg_7_inst : DFFR_X1 port map( D => n197, CK => clk, RN => n18, Q => 
                           IR_7_port, QN => n150);
   IR_reg_8_inst : DFFR_X1 port map( D => n198, CK => clk, RN => n18, Q => 
                           IR_8_port, QN => n149);
   IR_reg_9_inst : DFFR_X1 port map( D => n199, CK => clk, RN => n18, Q => 
                           IR_9_port, QN => n148);
   IR_reg_10_inst : DFFR_X1 port map( D => n200, CK => clk, RN => n18, Q => 
                           IR_10_port, QN => n147);
   IR_reg_11_inst : DFFR_X1 port map( D => n201, CK => clk, RN => n19, Q => 
                           IR_11_port, QN => n146);
   IR_reg_12_inst : DFFR_X1 port map( D => n202, CK => clk, RN => n19, Q => 
                           IR_12_port, QN => n145);
   IR_reg_13_inst : DFFR_X1 port map( D => n203, CK => clk, RN => n20, Q => 
                           IR_13_port, QN => n144);
   IR_reg_14_inst : DFFR_X1 port map( D => n204, CK => clk, RN => n20, Q => 
                           IR_14_port, QN => n143);
   IR_reg_15_inst : DFFR_X1 port map( D => n205, CK => clk, RN => n22, Q => 
                           IR_15_port, QN => n142);
   IR_reg_16_inst : DFFR_X1 port map( D => n206, CK => clk, RN => n22, Q => 
                           IR_16_port, QN => n141);
   IR_reg_17_inst : DFFR_X1 port map( D => n207, CK => clk, RN => n22, Q => 
                           IR_17_port, QN => n140);
   IR_reg_18_inst : DFFR_X1 port map( D => n208, CK => clk, RN => n22, Q => 
                           IR_18_port, QN => n139);
   IR_reg_19_inst : DFFR_X1 port map( D => n209, CK => clk, RN => n22, Q => 
                           IR_19_port, QN => n138);
   IR_reg_20_inst : DFFR_X1 port map( D => n210, CK => clk, RN => n23, Q => 
                           IR_20_port, QN => n137);
   IR_reg_21_inst : DFFR_X1 port map( D => n211, CK => clk, RN => n23, Q => 
                           IR_21_port, QN => n136);
   IR_reg_22_inst : DFFR_X1 port map( D => n212, CK => clk, RN => n23, Q => 
                           IR_22_port, QN => n135);
   IR_reg_23_inst : DFFR_X1 port map( D => n213, CK => clk, RN => n23, Q => 
                           IR_23_port, QN => n134);
   IR_reg_24_inst : DFFR_X1 port map( D => n214, CK => clk, RN => n23, Q => 
                           IR_24_port, QN => n133);
   IR_reg_25_inst : DFFR_X1 port map( D => n215, CK => clk, RN => n23, Q => 
                           IR_25_port, QN => n132);
   IR_reg_26_inst : DFFR_X1 port map( D => n216, CK => clk, RN => n23, Q => 
                           IR_26_port, QN => n131);
   IR_reg_27_inst : DFFR_X1 port map( D => n217, CK => clk, RN => n24, Q => 
                           IR_27_port, QN => n130);
   IR_reg_28_inst : DFFR_X1 port map( D => n218, CK => clk, RN => n24, Q => 
                           IR_28_port, QN => n129);
   IR_reg_29_inst : DFFR_X1 port map( D => n219, CK => clk, RN => n24, Q => 
                           IR_29_port, QN => n128);
   IR_reg_30_inst : DFFR_X1 port map( D => n220, CK => clk, RN => n24, Q => 
                           IR_30_port, QN => n127);
   IR_reg_31_inst : DFFR_X1 port map( D => n221, CK => clk, RN => n24, Q => 
                           IR_31_port, QN => n126);
   PCPlus4_reg_0_inst : DFFR_X1 port map( D => n189, CK => clk, RN => n16, Q =>
                           PCPlus4_0_port, QN => n125);
   PCPlus4_reg_1_inst : DFFR_X1 port map( D => n188, CK => clk, RN => n16, Q =>
                           PCPlus4_1_port, QN => n124);
   PCPlus4_reg_2_inst : DFFR_X1 port map( D => n187, CK => clk, RN => n16, Q =>
                           PCPlus4_2_port, QN => n123);
   PCPlus4_reg_3_inst : DFFR_X1 port map( D => n186, CK => clk, RN => n16, Q =>
                           PCPlus4_3_port, QN => n122);
   PCPlus4_reg_4_inst : DFFR_X1 port map( D => n185, CK => clk, RN => n16, Q =>
                           PCPlus4_4_port, QN => n121);
   PCPlus4_reg_5_inst : DFFR_X1 port map( D => n184, CK => clk, RN => n16, Q =>
                           PCPlus4_5_port, QN => n120);
   PCPlus4_reg_6_inst : DFFR_X1 port map( D => n183, CK => clk, RN => n16, Q =>
                           PCPlus4_6_port, QN => n119);
   PCPlus4_reg_7_inst : DFFR_X1 port map( D => n182, CK => clk, RN => n16, Q =>
                           PCPlus4_7_port, QN => n118);
   PCPlus4_reg_8_inst : DFFR_X1 port map( D => n181, CK => clk, RN => n16, Q =>
                           PCPlus4_8_port, QN => n117);
   PCPlus4_reg_9_inst : DFFR_X1 port map( D => n180, CK => clk, RN => n16, Q =>
                           PCPlus4_9_port, QN => n116);
   PCPlus4_reg_10_inst : DFFR_X1 port map( D => n179, CK => clk, RN => n16, Q 
                           => PCPlus4_10_port, QN => n115);
   PCPlus4_reg_11_inst : DFFR_X1 port map( D => n178, CK => clk, RN => n16, Q 
                           => PCPlus4_11_port, QN => n114);
   PCPlus4_reg_12_inst : DFFR_X1 port map( D => n177, CK => clk, RN => n15, Q 
                           => PCPlus4_12_port, QN => n113);
   PCPlus4_reg_13_inst : DFFR_X1 port map( D => n176, CK => clk, RN => n15, Q 
                           => PCPlus4_13_port, QN => n112);
   PCPlus4_reg_14_inst : DFFR_X1 port map( D => n175, CK => clk, RN => n15, Q 
                           => PCPlus4_14_port, QN => n111);
   PCPlus4_reg_15_inst : DFFR_X1 port map( D => n174, CK => clk, RN => n15, Q 
                           => PCPlus4_15_port, QN => n110);
   PCPlus4_reg_16_inst : DFFR_X1 port map( D => n173, CK => clk, RN => n15, Q 
                           => PCPlus4_16_port, QN => n109);
   PCPlus4_reg_17_inst : DFFR_X1 port map( D => n172, CK => clk, RN => n15, Q 
                           => PCPlus4_17_port, QN => n108);
   PCPlus4_reg_18_inst : DFFR_X1 port map( D => n171, CK => clk, RN => n15, Q 
                           => PCPlus4_18_port, QN => n107);
   PCPlus4_reg_19_inst : DFFR_X1 port map( D => n170, CK => clk, RN => n15, Q 
                           => PCPlus4_19_port, QN => n106);
   PCPlus4_reg_20_inst : DFFR_X1 port map( D => n169, CK => clk, RN => n15, Q 
                           => PCPlus4_20_port, QN => n105);
   PCPlus4_reg_21_inst : DFFR_X1 port map( D => n168, CK => clk, RN => n15, Q 
                           => PCPlus4_21_port, QN => n104);
   PCPlus4_reg_22_inst : DFFR_X1 port map( D => n167, CK => clk, RN => n15, Q 
                           => PCPlus4_22_port, QN => n103);
   PCPlus4_reg_23_inst : DFFR_X1 port map( D => n166, CK => clk, RN => n15, Q 
                           => PCPlus4_23_port, QN => n102);
   PCPlus4_reg_24_inst : DFFR_X1 port map( D => n165, CK => clk, RN => n14, Q 
                           => PCPlus4_24_port, QN => n101);
   PCPlus4_reg_25_inst : DFFR_X1 port map( D => n164, CK => clk, RN => n14, Q 
                           => PCPlus4_25_port, QN => n100);
   PCPlus4_reg_26_inst : DFFR_X1 port map( D => n163, CK => clk, RN => n14, Q 
                           => PCPlus4_26_port, QN => n99);
   PCPlus4_reg_27_inst : DFFR_X1 port map( D => n162, CK => clk, RN => n14, Q 
                           => PCPlus4_27_port, QN => n98);
   PCPlus4_reg_28_inst : DFFR_X1 port map( D => n161, CK => clk, RN => n14, Q 
                           => PCPlus4_28_port, QN => n97);
   PCPlus4_reg_29_inst : DFFR_X1 port map( D => n160, CK => clk, RN => n14, Q 
                           => PCPlus4_29_port, QN => n96);
   PCPlus4_reg_30_inst : DFFR_X1 port map( D => n159, CK => clk, RN => n14, Q 
                           => PCPlus4_30_port, QN => n95);
   PCPlus4_reg_31_inst : DFFR_X1 port map( D => n158, CK => clk, RN => n14, Q 
                           => PCPlus4_31_port, QN => n94);
   SignImmD_reg_0_inst : DFFR_X1 port map( D => SignImmD_wire_0_port, CK => clk
                           , RN => n17, Q => SignImmD_0_port, QN => n_1614);
   SignImmD_reg_1_inst : DFFR_X1 port map( D => SignImmD_wire_1_port, CK => clk
                           , RN => n17, Q => SignImmD_1_port, QN => n_1615);
   SignImmD_reg_2_inst : DFFR_X1 port map( D => SignImmD_wire_2_port, CK => clk
                           , RN => n17, Q => SignImmD_2_port, QN => n_1616);
   SignImmD_reg_3_inst : DFFR_X1 port map( D => SignImmD_wire_3_port, CK => clk
                           , RN => n17, Q => SignImmD_3_port, QN => n_1617);
   SignImmD_reg_4_inst : DFFR_X1 port map( D => SignImmD_wire_4_port, CK => clk
                           , RN => n17, Q => SignImmD_4_port, QN => n_1618);
   SignImmD_reg_5_inst : DFFR_X1 port map( D => SignImmD_wire_5_port, CK => clk
                           , RN => n17, Q => SignImmD_5_port, QN => n_1619);
   SignImmD_reg_6_inst : DFFR_X1 port map( D => SignImmD_wire_6_port, CK => clk
                           , RN => n18, Q => SignImmD_6_port, QN => n_1620);
   SignImmD_reg_7_inst : DFFR_X1 port map( D => SignImmD_wire_7_port, CK => clk
                           , RN => n18, Q => SignImmD_7_port, QN => n_1621);
   SignImmD_reg_8_inst : DFFR_X1 port map( D => SignImmD_wire_8_port, CK => clk
                           , RN => n18, Q => SignImmD_8_port, QN => n_1622);
   SignImmD_reg_9_inst : DFFR_X1 port map( D => SignImmD_wire_9_port, CK => clk
                           , RN => n18, Q => SignImmD_9_port, QN => n_1623);
   SignImmD_reg_10_inst : DFFR_X1 port map( D => SignImmD_wire_10_port, CK => 
                           clk, RN => n18, Q => SignImmD_10_port, QN => n_1624)
                           ;
   SignImmD_reg_11_inst : DFFR_X1 port map( D => SignImmD_wire_11_port, CK => 
                           clk, RN => n19, Q => SignImmD_11_port, QN => n_1625)
                           ;
   SignImmD_reg_12_inst : DFFR_X1 port map( D => SignImmD_wire_12_port, CK => 
                           clk, RN => n19, Q => SignImmD_12_port, QN => n_1626)
                           ;
   SignImmD_reg_13_inst : DFFR_X1 port map( D => SignImmD_wire_13_port, CK => 
                           clk, RN => n19, Q => SignImmD_13_port, QN => n_1627)
                           ;
   SignImmD_reg_14_inst : DFFR_X1 port map( D => SignImmD_wire_14_port, CK => 
                           clk, RN => n20, Q => SignImmD_14_port, QN => n_1628)
                           ;
   SignImmD_reg_15_inst : DFFR_X1 port map( D => SignImmD_wire_15_port, CK => 
                           clk, RN => n22, Q => SignImmD_15_port, QN => n_1629)
                           ;
   SignImmD_reg_16_inst : DFFR_X1 port map( D => SignImmD_wire_16_port, CK => 
                           clk, RN => n22, Q => SignImmD_16_port, QN => n_1630)
                           ;
   SignImmD_reg_17_inst : DFFR_X1 port map( D => SignImmD_wire_17_port, CK => 
                           clk, RN => n21, Q => SignImmD_17_port, QN => n_1631)
                           ;
   SignImmD_reg_18_inst : DFFR_X1 port map( D => SignImmD_wire_18_port, CK => 
                           clk, RN => n21, Q => SignImmD_18_port, QN => n_1632)
                           ;
   SignImmD_reg_19_inst : DFFR_X1 port map( D => SignImmD_wire_19_port, CK => 
                           clk, RN => n21, Q => SignImmD_19_port, QN => n_1633)
                           ;
   SignImmD_reg_20_inst : DFFR_X1 port map( D => SignImmD_wire_20_port, CK => 
                           clk, RN => n21, Q => SignImmD_20_port, QN => n_1634)
                           ;
   SignImmD_reg_21_inst : DFFR_X1 port map( D => SignImmD_wire_21_port, CK => 
                           clk, RN => n21, Q => SignImmD_21_port, QN => n_1635)
                           ;
   SignImmD_reg_22_inst : DFFR_X1 port map( D => SignImmD_wire_22_port, CK => 
                           clk, RN => n21, Q => SignImmD_22_port, QN => n_1636)
                           ;
   SignImmD_reg_23_inst : DFFR_X1 port map( D => SignImmD_wire_23_port, CK => 
                           clk, RN => n21, Q => SignImmD_23_port, QN => n_1637)
                           ;
   SignImmD_reg_24_inst : DFFR_X1 port map( D => SignImmD_wire_24_port, CK => 
                           clk, RN => n21, Q => SignImmD_24_port, QN => n_1638)
                           ;
   SignImmD_reg_25_inst : DFFR_X1 port map( D => SignImmD_wire_25_port, CK => 
                           clk, RN => n21, Q => SignImmD_25_port, QN => n_1639)
                           ;
   SignImmD_reg_26_inst : DFFR_X1 port map( D => SignImmD_wire_26_port, CK => 
                           clk, RN => n21, Q => SignImmD_26_port, QN => n_1640)
                           ;
   SignImmD_reg_27_inst : DFFR_X1 port map( D => SignImmD_wire_27_port, CK => 
                           clk, RN => n21, Q => SignImmD_27_port, QN => n_1641)
                           ;
   SignImmD_reg_28_inst : DFFR_X1 port map( D => SignImmD_wire_28_port, CK => 
                           clk, RN => n21, Q => SignImmD_28_port, QN => n_1642)
                           ;
   SignImmD_reg_29_inst : DFFR_X1 port map( D => SignImmD_wire_29_port, CK => 
                           clk, RN => n20, Q => SignImmD_29_port, QN => n_1643)
                           ;
   SignImmD_reg_30_inst : DFFR_X1 port map( D => SignImmD_wire_30_port, CK => 
                           clk, RN => n20, Q => SignImmD_30_port, QN => n_1644)
                           ;
   SignImmD_reg_31_inst : DFFR_X1 port map( D => SignImmD_wire_31_port, CK => 
                           clk, RN => n20, Q => SignImmD_31_port, QN => n_1645)
                           ;
   RdD_reg_0_inst : DFFR_X1 port map( D => RdD_wire_0_port, CK => clk, RN => 
                           n19, Q => RdD_0_port, QN => n_1646);
   RdD_reg_1_inst : DFFR_X1 port map( D => RdD_wire_1_port, CK => clk, RN => 
                           n19, Q => RdD_1_port, QN => n_1647);
   RdD_reg_2_inst : DFFR_X1 port map( D => RdD_wire_2_port, CK => clk, RN => 
                           n19, Q => RdD_2_port, QN => n_1648);
   RdD_reg_3_inst : DFFR_X1 port map( D => RdD_wire_3_port, CK => clk, RN => 
                           n20, Q => RdD_3_port, QN => n_1649);
   RdD_reg_4_inst : DFFR_X1 port map( D => RdD_wire_4_port, CK => clk, RN => 
                           n20, Q => RdD_4_port, QN => n_1650);
   RtD_reg_0_inst : DFFR_X1 port map( D => RtD_H_0_port, CK => clk, RN => n22, 
                           Q => RtD_0_port, QN => n_1651);
   RtD_reg_1_inst : DFFR_X1 port map( D => RtD_H_1_port, CK => clk, RN => n22, 
                           Q => RtD_1_port, QN => n_1652);
   RtD_reg_2_inst : DFFR_X1 port map( D => RtD_H_2_port, CK => clk, RN => n22, 
                           Q => RtD_2_port, QN => n_1653);
   RtD_reg_3_inst : DFFR_X1 port map( D => RtD_H_3_port, CK => clk, RN => n22, 
                           Q => RtD_3_port, QN => n_1654);
   RtD_reg_4_inst : DFFR_X1 port map( D => RtD_H_4_port, CK => clk, RN => n22, 
                           Q => RtD_4_port, QN => n_1655);
   RsD_reg_0_inst : DFFR_X1 port map( D => RsD_H_0_port, CK => clk, RN => n23, 
                           Q => RsD_0_port, QN => n_1656);
   RsD_reg_1_inst : DFFR_X1 port map( D => RsD_H_1_port, CK => clk, RN => n23, 
                           Q => RsD_1_port, QN => n_1657);
   RsD_reg_2_inst : DFFR_X1 port map( D => RsD_H_2_port, CK => clk, RN => n23, 
                           Q => RsD_2_port, QN => n_1658);
   RsD_reg_3_inst : DFFR_X1 port map( D => RsD_H_3_port, CK => clk, RN => n23, 
                           Q => RsD_3_port, QN => n_1659);
   RsD_reg_4_inst : DFFR_X1 port map( D => RsD_H_4_port, CK => clk, RN => n23, 
                           Q => RsD_4_port, QN => n_1660);
   WriteDataE_reg_0_inst : DFFR_X1 port map( D => WriteDataE_wire_0_port, CK =>
                           clk, RN => n1, Q => WriteDataE_0_port, QN => n_1661)
                           ;
   WriteDataE_reg_1_inst : DFFR_X1 port map( D => WriteDataE_wire_1_port, CK =>
                           clk, RN => n1, Q => WriteDataE_1_port, QN => n_1662)
                           ;
   WriteDataE_reg_2_inst : DFFR_X1 port map( D => WriteDataE_wire_2_port, CK =>
                           clk, RN => n1, Q => WriteDataE_2_port, QN => n_1663)
                           ;
   WriteDataE_reg_3_inst : DFFR_X1 port map( D => WriteDataE_wire_3_port, CK =>
                           clk, RN => n2, Q => WriteDataE_3_port, QN => n_1664)
                           ;
   WriteDataE_reg_4_inst : DFFR_X1 port map( D => WriteDataE_wire_4_port, CK =>
                           clk, RN => n13, Q => WriteDataE_4_port, QN => n_1665
                           );
   WriteDataE_reg_5_inst : DFFR_X1 port map( D => WriteDataE_wire_5_port, CK =>
                           clk, RN => n5, Q => WriteDataE_5_port, QN => n_1666)
                           ;
   WriteDataE_reg_6_inst : DFFR_X1 port map( D => WriteDataE_wire_6_port, CK =>
                           clk, RN => n2, Q => WriteDataE_6_port, QN => n_1667)
                           ;
   WriteDataE_reg_7_inst : DFFR_X1 port map( D => WriteDataE_wire_7_port, CK =>
                           clk, RN => n2, Q => WriteDataE_7_port, QN => n_1668)
                           ;
   WriteDataE_reg_8_inst : DFFR_X1 port map( D => WriteDataE_wire_8_port, CK =>
                           clk, RN => n4, Q => WriteDataE_8_port, QN => n_1669)
                           ;
   WriteDataE_reg_9_inst : DFFR_X1 port map( D => WriteDataE_wire_9_port, CK =>
                           clk, RN => n12, Q => WriteDataE_9_port, QN => n_1670
                           );
   WriteDataE_reg_10_inst : DFFR_X1 port map( D => WriteDataE_wire_10_port, CK 
                           => clk, RN => n3, Q => WriteDataE_10_port, QN => 
                           n_1671);
   WriteDataE_reg_11_inst : DFFR_X1 port map( D => WriteDataE_wire_11_port, CK 
                           => clk, RN => n4, Q => WriteDataE_11_port, QN => 
                           n_1672);
   WriteDataE_reg_12_inst : DFFR_X1 port map( D => WriteDataE_wire_12_port, CK 
                           => clk, RN => n11, Q => WriteDataE_12_port, QN => 
                           n_1673);
   WriteDataE_reg_13_inst : DFFR_X1 port map( D => WriteDataE_wire_13_port, CK 
                           => clk, RN => n3, Q => WriteDataE_13_port, QN => 
                           n_1674);
   WriteDataE_reg_14_inst : DFFR_X1 port map( D => WriteDataE_wire_14_port, CK 
                           => clk, RN => n4, Q => WriteDataE_14_port, QN => 
                           n_1675);
   WriteDataE_reg_15_inst : DFFR_X1 port map( D => WriteDataE_wire_15_port, CK 
                           => clk, RN => n6, Q => WriteDataE_15_port, QN => 
                           n_1676);
   WriteDataE_reg_16_inst : DFFR_X1 port map( D => WriteDataE_wire_16_port, CK 
                           => clk, RN => n13, Q => WriteDataE_16_port, QN => 
                           n_1677);
   WriteDataE_reg_17_inst : DFFR_X1 port map( D => WriteDataE_wire_17_port, CK 
                           => clk, RN => n7, Q => WriteDataE_17_port, QN => 
                           n_1678);
   WriteDataE_reg_18_inst : DFFR_X1 port map( D => WriteDataE_wire_18_port, CK 
                           => clk, RN => n7, Q => WriteDataE_18_port, QN => 
                           n_1679);
   WriteDataE_reg_19_inst : DFFR_X1 port map( D => WriteDataE_wire_19_port, CK 
                           => clk, RN => n7, Q => WriteDataE_19_port, QN => 
                           n_1680);
   WriteDataE_reg_20_inst : DFFR_X1 port map( D => WriteDataE_wire_20_port, CK 
                           => clk, RN => n8, Q => WriteDataE_20_port, QN => 
                           n_1681);
   WriteDataE_reg_21_inst : DFFR_X1 port map( D => WriteDataE_wire_21_port, CK 
                           => clk, RN => n8, Q => WriteDataE_21_port, QN => 
                           n_1682);
   WriteDataE_reg_22_inst : DFFR_X1 port map( D => WriteDataE_wire_22_port, CK 
                           => clk, RN => n9, Q => WriteDataE_22_port, QN => 
                           n_1683);
   WriteDataE_reg_23_inst : DFFR_X1 port map( D => WriteDataE_wire_23_port, CK 
                           => clk, RN => n9, Q => WriteDataE_23_port, QN => 
                           n_1684);
   WriteDataE_reg_24_inst : DFFR_X1 port map( D => WriteDataE_wire_24_port, CK 
                           => clk, RN => n11, Q => WriteDataE_24_port, QN => 
                           n_1685);
   WriteDataE_reg_25_inst : DFFR_X1 port map( D => WriteDataE_wire_25_port, CK 
                           => clk, RN => n9, Q => WriteDataE_25_port, QN => 
                           n_1686);
   WriteDataE_reg_26_inst : DFFR_X1 port map( D => WriteDataE_wire_26_port, CK 
                           => clk, RN => n10, Q => WriteDataE_26_port, QN => 
                           n_1687);
   WriteDataE_reg_27_inst : DFFR_X1 port map( D => WriteDataE_wire_27_port, CK 
                           => clk, RN => n10, Q => WriteDataE_27_port, QN => 
                           n_1688);
   WriteDataE_reg_28_inst : DFFR_X1 port map( D => WriteDataE_wire_28_port, CK 
                           => clk, RN => n12, Q => WriteDataE_28_port, QN => 
                           n_1689);
   WriteDataE_reg_29_inst : DFFR_X1 port map( D => WriteDataE_wire_29_port, CK 
                           => clk, RN => n5, Q => WriteDataE_29_port, QN => 
                           n_1690);
   WriteDataE_reg_30_inst : DFFR_X1 port map( D => WriteDataE_wire_30_port, CK 
                           => clk, RN => n6, Q => WriteDataE_30_port, QN => 
                           n_1691);
   WriteDataE_reg_31_inst : DFFR_X1 port map( D => WriteDataE_wire_31_port, CK 
                           => clk, RN => n12, Q => WriteDataE_31_port, QN => 
                           n_1692);
   WriteRegE_reg_0_inst : DFFR_X1 port map( D => WriteRegE_H_0_port, CK => clk,
                           RN => n18, Q => WriteRegE_0_port, QN => n_1693);
   WriteRegE_reg_1_inst : DFFR_X1 port map( D => WriteRegE_H_1_port, CK => clk,
                           RN => n19, Q => WriteRegE_1_port, QN => n_1694);
   WriteRegE_reg_2_inst : DFFR_X1 port map( D => WriteRegE_H_2_port, CK => clk,
                           RN => n19, Q => WriteRegE_2_port, QN => n_1695);
   WriteRegE_reg_3_inst : DFFR_X1 port map( D => WriteRegE_H_3_port, CK => clk,
                           RN => n20, Q => WriteRegE_3_port, QN => n_1696);
   WriteRegE_reg_4_inst : DFFR_X1 port map( D => WriteRegE_H_4_port, CK => clk,
                           RN => n20, Q => WriteRegE_4_port, QN => n_1697);
   ALUOutE_reg_0_inst : DFFR_X1 port map( D => ALUOutE_wire_0_port, CK => clk, 
                           RN => n14, Q => ALUOutE_0_port, QN => n_1698);
   ALUOutE_reg_1_inst : DFFR_X1 port map( D => ALUOutE_wire_1_port, CK => clk, 
                           RN => n1, Q => ALUOutE_1_port, QN => n_1699);
   ALUOutE_reg_2_inst : DFFR_X1 port map( D => ALUOutE_wire_2_port, CK => clk, 
                           RN => n1, Q => ALUOutE_2_port, QN => n_1700);
   ALUOutE_reg_3_inst : DFFR_X1 port map( D => ALUOutE_wire_3_port, CK => clk, 
                           RN => n2, Q => ALUOutE_3_port, QN => n_1701);
   ALUOutE_reg_4_inst : DFFR_X1 port map( D => ALUOutE_wire_4_port, CK => clk, 
                           RN => n13, Q => ALUOutE_4_port, QN => n_1702);
   ALUOutE_reg_5_inst : DFFR_X1 port map( D => ALUOutE_wire_5_port, CK => clk, 
                           RN => n5, Q => ALUOutE_5_port, QN => n_1703);
   ALUOutE_reg_6_inst : DFFR_X1 port map( D => ALUOutE_wire_6_port, CK => clk, 
                           RN => n2, Q => ALUOutE_6_port, QN => n_1704);
   ALUOutE_reg_7_inst : DFFR_X1 port map( D => ALUOutE_wire_7_port, CK => clk, 
                           RN => n3, Q => ALUOutE_7_port, QN => n_1705);
   ALUOutE_reg_8_inst : DFFR_X1 port map( D => ALUOutE_wire_8_port, CK => clk, 
                           RN => n5, Q => ALUOutE_8_port, QN => n_1706);
   ALUOutE_reg_9_inst : DFFR_X1 port map( D => ALUOutE_wire_9_port, CK => clk, 
                           RN => n12, Q => ALUOutE_9_port, QN => n_1707);
   ALUOutE_reg_10_inst : DFFR_X1 port map( D => ALUOutE_wire_10_port, CK => clk
                           , RN => n3, Q => ALUOutE_10_port, QN => n_1708);
   ALUOutE_reg_11_inst : DFFR_X1 port map( D => ALUOutE_wire_11_port, CK => clk
                           , RN => n4, Q => ALUOutE_11_port, QN => n_1709);
   ALUOutE_reg_12_inst : DFFR_X1 port map( D => ALUOutE_wire_12_port, CK => clk
                           , RN => n11, Q => ALUOutE_12_port, QN => n_1710);
   ALUOutE_reg_13_inst : DFFR_X1 port map( D => ALUOutE_wire_13_port, CK => clk
                           , RN => n3, Q => ALUOutE_13_port, QN => n_1711);
   ALUOutE_reg_14_inst : DFFR_X1 port map( D => ALUOutE_wire_14_port, CK => clk
                           , RN => n4, Q => ALUOutE_14_port, QN => n_1712);
   ALUOutE_reg_15_inst : DFFR_X1 port map( D => ALUOutE_wire_15_port, CK => clk
                           , RN => n6, Q => ALUOutE_15_port, QN => n_1713);
   ALUOutE_reg_16_inst : DFFR_X1 port map( D => ALUOutE_wire_16_port, CK => clk
                           , RN => n13, Q => ALUOutE_16_port, QN => n_1714);
   ALUOutE_reg_17_inst : DFFR_X1 port map( D => ALUOutE_wire_17_port, CK => clk
                           , RN => n7, Q => ALUOutE_17_port, QN => n_1715);
   ALUOutE_reg_18_inst : DFFR_X1 port map( D => ALUOutE_wire_18_port, CK => clk
                           , RN => n7, Q => ALUOutE_18_port, QN => n_1716);
   ALUOutE_reg_19_inst : DFFR_X1 port map( D => ALUOutE_wire_19_port, CK => clk
                           , RN => n8, Q => ALUOutE_19_port, QN => n_1717);
   ALUOutE_reg_20_inst : DFFR_X1 port map( D => ALUOutE_wire_20_port, CK => clk
                           , RN => n8, Q => ALUOutE_20_port, QN => n_1718);
   ALUOutE_reg_21_inst : DFFR_X1 port map( D => ALUOutE_wire_21_port, CK => clk
                           , RN => n8, Q => ALUOutE_21_port, QN => n_1719);
   ALUOutE_reg_22_inst : DFFR_X1 port map( D => ALUOutE_wire_22_port, CK => clk
                           , RN => n9, Q => ALUOutE_22_port, QN => n_1720);
   ALUOutE_reg_23_inst : DFFR_X1 port map( D => ALUOutE_wire_23_port, CK => clk
                           , RN => n9, Q => ALUOutE_23_port, QN => n_1721);
   ALUOutE_reg_24_inst : DFFR_X1 port map( D => ALUOutE_wire_24_port, CK => clk
                           , RN => n11, Q => ALUOutE_24_port, QN => n_1722);
   ALUOutE_reg_25_inst : DFFR_X1 port map( D => ALUOutE_wire_25_port, CK => clk
                           , RN => n10, Q => ALUOutE_25_port, QN => n_1723);
   ALUOutE_reg_26_inst : DFFR_X1 port map( D => ALUOutE_wire_26_port, CK => clk
                           , RN => n10, Q => ALUOutE_26_port, QN => n_1724);
   ALUOutE_reg_27_inst : DFFR_X1 port map( D => ALUOutE_wire_27_port, CK => clk
                           , RN => n11, Q => ALUOutE_27_port, QN => n_1725);
   ALUOutE_reg_28_inst : DFFR_X1 port map( D => ALUOutE_wire_28_port, CK => clk
                           , RN => n13, Q => ALUOutE_28_port, QN => n_1726);
   ALUOutE_reg_29_inst : DFFR_X1 port map( D => ALUOutE_wire_29_port, CK => clk
                           , RN => n6, Q => ALUOutE_29_port, QN => n_1727);
   ALUOutE_reg_30_inst : DFFR_X1 port map( D => ALUOutE_wire_30_port, CK => clk
                           , RN => n6, Q => ALUOutE_30_port, QN => n_1728);
   ALUOutE_reg_31_inst : DFFR_X1 port map( D => ALUOutE_wire_31_port, CK => clk
                           , RN => n12, Q => ALUOutE_31_port, QN => n_1729);
   WriteRegM_reg_0_inst : DFFR_X1 port map( D => WriteRegMOut_H_0_port, CK => 
                           clk, RN => n18, Q => WriteRegM_0_port, QN => n_1730)
                           ;
   WriteRegM_reg_1_inst : DFFR_X1 port map( D => WriteRegMOut_H_1_port, CK => 
                           clk, RN => n19, Q => WriteRegM_1_port, QN => n_1731)
                           ;
   WriteRegM_reg_2_inst : DFFR_X1 port map( D => WriteRegMOut_H_2_port, CK => 
                           clk, RN => n19, Q => WriteRegM_2_port, QN => n_1732)
                           ;
   WriteRegM_reg_3_inst : DFFR_X1 port map( D => WriteRegMOut_H_3_port, CK => 
                           clk, RN => n20, Q => WriteRegM_3_port, QN => n_1733)
                           ;
   WriteRegM_reg_4_inst : DFFR_X1 port map( D => WriteRegMOut_H_4_port, CK => 
                           clk, RN => n20, Q => WriteRegM_4_port, QN => n_1734)
                           ;
   ALUOutM_reg_1_inst : DFFR_X1 port map( D => ALUOutMOut_wire_1_port, CK => 
                           clk, RN => n1, Q => ALUOutM_1_port, QN => n_1735);
   ALUOutM_reg_2_inst : DFFR_X1 port map( D => ALUOutMOut_wire_2_port, CK => 
                           clk, RN => n1, Q => ALUOutM_2_port, QN => n_1736);
   ALUOutM_reg_3_inst : DFFR_X1 port map( D => ALUOutMOut_wire_3_port, CK => 
                           clk, RN => n2, Q => ALUOutM_3_port, QN => n_1737);
   ALUOutM_reg_4_inst : DFFR_X1 port map( D => ALUOutMOut_wire_4_port, CK => 
                           clk, RN => n13, Q => ALUOutM_4_port, QN => n_1738);
   ALUOutM_reg_5_inst : DFFR_X1 port map( D => ALUOutMOut_wire_5_port, CK => 
                           clk, RN => n5, Q => ALUOutM_5_port, QN => n_1739);
   ALUOutM_reg_6_inst : DFFR_X1 port map( D => ALUOutMOut_wire_6_port, CK => 
                           clk, RN => n2, Q => ALUOutM_6_port, QN => n_1740);
   ALUOutM_reg_7_inst : DFFR_X1 port map( D => ALUOutMOut_wire_7_port, CK => 
                           clk, RN => n3, Q => ALUOutM_7_port, QN => n_1741);
   ALUOutM_reg_8_inst : DFFR_X1 port map( D => ALUOutMOut_wire_8_port, CK => 
                           clk, RN => n5, Q => ALUOutM_8_port, QN => n_1742);
   ALUOutM_reg_9_inst : DFFR_X1 port map( D => ALUOutMOut_wire_9_port, CK => 
                           clk, RN => n12, Q => ALUOutM_9_port, QN => n_1743);
   ALUOutM_reg_10_inst : DFFR_X1 port map( D => ALUOutMOut_wire_10_port, CK => 
                           clk, RN => n3, Q => ALUOutM_10_port, QN => n_1744);
   ALUOutM_reg_11_inst : DFFR_X1 port map( D => ALUOutMOut_wire_11_port, CK => 
                           clk, RN => n4, Q => ALUOutM_11_port, QN => n_1745);
   ALUOutM_reg_12_inst : DFFR_X1 port map( D => ALUOutMOut_wire_12_port, CK => 
                           clk, RN => n11, Q => ALUOutM_12_port, QN => n_1746);
   ALUOutM_reg_13_inst : DFFR_X1 port map( D => ALUOutMOut_wire_13_port, CK => 
                           clk, RN => n3, Q => ALUOutM_13_port, QN => n_1747);
   ALUOutM_reg_14_inst : DFFR_X1 port map( D => ALUOutMOut_wire_14_port, CK => 
                           clk, RN => n4, Q => ALUOutM_14_port, QN => n_1748);
   ALUOutM_reg_15_inst : DFFR_X1 port map( D => ALUOutMOut_wire_15_port, CK => 
                           clk, RN => n6, Q => ALUOutM_15_port, QN => n_1749);
   ALUOutM_reg_16_inst : DFFR_X1 port map( D => ALUOutMOut_wire_16_port, CK => 
                           clk, RN => n13, Q => ALUOutM_16_port, QN => n_1750);
   ALUOutM_reg_17_inst : DFFR_X1 port map( D => ALUOutMOut_wire_17_port, CK => 
                           clk, RN => n7, Q => ALUOutM_17_port, QN => n_1751);
   ALUOutM_reg_18_inst : DFFR_X1 port map( D => ALUOutMOut_wire_18_port, CK => 
                           clk, RN => n7, Q => ALUOutM_18_port, QN => n_1752);
   ALUOutM_reg_19_inst : DFFR_X1 port map( D => ALUOutMOut_wire_19_port, CK => 
                           clk, RN => n8, Q => ALUOutM_19_port, QN => n_1753);
   ALUOutM_reg_20_inst : DFFR_X1 port map( D => ALUOutMOut_wire_20_port, CK => 
                           clk, RN => n8, Q => ALUOutM_20_port, QN => n_1754);
   ALUOutM_reg_21_inst : DFFR_X1 port map( D => ALUOutMOut_wire_21_port, CK => 
                           clk, RN => n8, Q => ALUOutM_21_port, QN => n_1755);
   ALUOutM_reg_22_inst : DFFR_X1 port map( D => ALUOutMOut_wire_22_port, CK => 
                           clk, RN => n9, Q => ALUOutM_22_port, QN => n_1756);
   ALUOutM_reg_23_inst : DFFR_X1 port map( D => ALUOutMOut_wire_23_port, CK => 
                           clk, RN => n9, Q => ALUOutM_23_port, QN => n_1757);
   ALUOutM_reg_24_inst : DFFR_X1 port map( D => ALUOutMOut_wire_24_port, CK => 
                           clk, RN => n11, Q => ALUOutM_24_port, QN => n_1758);
   ALUOutM_reg_25_inst : DFFR_X1 port map( D => ALUOutMOut_wire_25_port, CK => 
                           clk, RN => n10, Q => ALUOutM_25_port, QN => n_1759);
   ALUOutM_reg_26_inst : DFFR_X1 port map( D => ALUOutMOut_wire_26_port, CK => 
                           clk, RN => n10, Q => ALUOutM_26_port, QN => n_1760);
   ALUOutM_reg_27_inst : DFFR_X1 port map( D => ALUOutMOut_wire_27_port, CK => 
                           clk, RN => n10, Q => ALUOutM_27_port, QN => n_1761);
   ALUOutM_reg_28_inst : DFFR_X1 port map( D => ALUOutMOut_wire_28_port, CK => 
                           clk, RN => n13, Q => ALUOutM_28_port, QN => n_1762);
   ALUOutM_reg_29_inst : DFFR_X1 port map( D => ALUOutMOut_wire_29_port, CK => 
                           clk, RN => n5, Q => ALUOutM_29_port, QN => n_1763);
   ALUOutM_reg_30_inst : DFFR_X1 port map( D => ALUOutMOut_wire_30_port, CK => 
                           clk, RN => n6, Q => ALUOutM_30_port, QN => n_1764);
   ALUOutM_reg_31_inst : DFFR_X1 port map( D => ALUOutMOut_wire_31_port, CK => 
                           clk, RN => n12, Q => ALUOutM_31_port, QN => n_1765);
   ReadDataM_reg_0_inst : DFFR_X1 port map( D => ReadDataM_wire_0_port, CK => 
                           clk, RN => n24, Q => ReadDataM_0_port, QN => n_1766)
                           ;
   ReadDataM_reg_1_inst : DFFR_X1 port map( D => ReadDataM_wire_1_port, CK => 
                           clk, RN => n24, Q => ReadDataM_1_port, QN => n_1767)
                           ;
   ReadDataM_reg_2_inst : DFFR_X1 port map( D => ReadDataM_wire_2_port, CK => 
                           clk, RN => n24, Q => ReadDataM_2_port, QN => n_1768)
                           ;
   ReadDataM_reg_3_inst : DFFR_X1 port map( D => ReadDataM_wire_3_port, CK => 
                           clk, RN => n24, Q => ReadDataM_3_port, QN => n_1769)
                           ;
   ReadDataM_reg_4_inst : DFFR_X1 port map( D => ReadDataM_wire_4_port, CK => 
                           clk, RN => n24, Q => ReadDataM_4_port, QN => n_1770)
                           ;
   ReadDataM_reg_5_inst : DFFR_X1 port map( D => ReadDataM_wire_5_port, CK => 
                           clk, RN => n24, Q => ReadDataM_5_port, QN => n_1771)
                           ;
   ReadDataM_reg_6_inst : DFFR_X1 port map( D => ReadDataM_wire_6_port, CK => 
                           clk, RN => n24, Q => ReadDataM_6_port, QN => n_1772)
                           ;
   ReadDataM_reg_7_inst : DFFR_X1 port map( D => ReadDataM_wire_7_port, CK => 
                           clk, RN => n25, Q => ReadDataM_7_port, QN => n_1773)
                           ;
   ReadDataM_reg_8_inst : DFFR_X1 port map( D => ReadDataM_wire_8_port, CK => 
                           clk, RN => n25, Q => ReadDataM_8_port, QN => n_1774)
                           ;
   ReadDataM_reg_9_inst : DFFR_X1 port map( D => ReadDataM_wire_9_port, CK => 
                           clk, RN => n25, Q => ReadDataM_9_port, QN => n_1775)
                           ;
   ReadDataM_reg_10_inst : DFFR_X1 port map( D => ReadDataM_wire_10_port, CK =>
                           clk, RN => n25, Q => ReadDataM_10_port, QN => n_1776
                           );
   ReadDataM_reg_11_inst : DFFR_X1 port map( D => ReadDataM_wire_11_port, CK =>
                           clk, RN => n25, Q => ReadDataM_11_port, QN => n_1777
                           );
   ReadDataM_reg_12_inst : DFFR_X1 port map( D => ReadDataM_wire_12_port, CK =>
                           clk, RN => n25, Q => ReadDataM_12_port, QN => n_1778
                           );
   ReadDataM_reg_13_inst : DFFR_X1 port map( D => ReadDataM_wire_13_port, CK =>
                           clk, RN => n25, Q => ReadDataM_13_port, QN => n_1779
                           );
   ReadDataM_reg_14_inst : DFFR_X1 port map( D => ReadDataM_wire_14_port, CK =>
                           clk, RN => n25, Q => ReadDataM_14_port, QN => n_1780
                           );
   ReadDataM_reg_15_inst : DFFR_X1 port map( D => ReadDataM_wire_15_port, CK =>
                           clk, RN => n25, Q => ReadDataM_15_port, QN => n_1781
                           );
   ReadDataM_reg_16_inst : DFFR_X1 port map( D => ReadDataM_wire_16_port, CK =>
                           clk, RN => n25, Q => ReadDataM_16_port, QN => n_1782
                           );
   ReadDataM_reg_17_inst : DFFR_X1 port map( D => ReadDataM_wire_17_port, CK =>
                           clk, RN => n25, Q => ReadDataM_17_port, QN => n_1783
                           );
   ReadDataM_reg_18_inst : DFFR_X1 port map( D => ReadDataM_wire_18_port, CK =>
                           clk, RN => n25, Q => ReadDataM_18_port, QN => n_1784
                           );
   ReadDataM_reg_19_inst : DFFR_X1 port map( D => ReadDataM_wire_19_port, CK =>
                           clk, RN => n26, Q => ReadDataM_19_port, QN => n_1785
                           );
   ReadDataM_reg_20_inst : DFFR_X1 port map( D => ReadDataM_wire_20_port, CK =>
                           clk, RN => n26, Q => ReadDataM_20_port, QN => n_1786
                           );
   ReadDataM_reg_21_inst : DFFR_X1 port map( D => ReadDataM_wire_21_port, CK =>
                           clk, RN => n26, Q => ReadDataM_21_port, QN => n_1787
                           );
   ReadDataM_reg_22_inst : DFFR_X1 port map( D => ReadDataM_wire_22_port, CK =>
                           clk, RN => n26, Q => ReadDataM_22_port, QN => n_1788
                           );
   ReadDataM_reg_23_inst : DFFR_X1 port map( D => ReadDataM_wire_23_port, CK =>
                           clk, RN => n26, Q => ReadDataM_23_port, QN => n_1789
                           );
   ReadDataM_reg_24_inst : DFFR_X1 port map( D => ReadDataM_wire_24_port, CK =>
                           clk, RN => n26, Q => ReadDataM_24_port, QN => n_1790
                           );
   ReadDataM_reg_25_inst : DFFR_X1 port map( D => ReadDataM_wire_25_port, CK =>
                           clk, RN => n26, Q => ReadDataM_25_port, QN => n_1791
                           );
   ReadDataM_reg_26_inst : DFFR_X1 port map( D => ReadDataM_wire_26_port, CK =>
                           clk, RN => n26, Q => ReadDataM_26_port, QN => n_1792
                           );
   ReadDataM_reg_27_inst : DFFR_X1 port map( D => ReadDataM_wire_27_port, CK =>
                           clk, RN => n26, Q => ReadDataM_27_port, QN => n_1793
                           );
   ReadDataM_reg_28_inst : DFFR_X1 port map( D => ReadDataM_wire_28_port, CK =>
                           clk, RN => n26, Q => ReadDataM_28_port, QN => n_1794
                           );
   ReadDataM_reg_29_inst : DFFR_X1 port map( D => ReadDataM_wire_29_port, CK =>
                           clk, RN => n26, Q => ReadDataM_29_port, QN => n_1795
                           );
   ReadDataM_reg_30_inst : DFFR_X1 port map( D => ReadDataM_wire_30_port, CK =>
                           clk, RN => n26, Q => ReadDataM_30_port, QN => n_1796
                           );
   ReadDataM_reg_31_inst : DFFR_X1 port map( D => ReadDataM_wire_31_port, CK =>
                           clk, RN => n222, Q => ReadDataM_31_port, QN => 
                           n_1797);
   fetch_stage : fetch_stage_wrapper_nbit32_nwords64 port map( PCBranchD(31) =>
                           PCBranchD_wire_31_port, PCBranchD(30) => 
                           PCBranchD_wire_30_port, PCBranchD(29) => 
                           PCBranchD_wire_29_port, PCBranchD(28) => 
                           PCBranchD_wire_28_port, PCBranchD(27) => 
                           PCBranchD_wire_27_port, PCBranchD(26) => 
                           PCBranchD_wire_26_port, PCBranchD(25) => 
                           PCBranchD_wire_25_port, PCBranchD(24) => 
                           PCBranchD_wire_24_port, PCBranchD(23) => 
                           PCBranchD_wire_23_port, PCBranchD(22) => 
                           PCBranchD_wire_22_port, PCBranchD(21) => 
                           PCBranchD_wire_21_port, PCBranchD(20) => 
                           PCBranchD_wire_20_port, PCBranchD(19) => 
                           PCBranchD_wire_19_port, PCBranchD(18) => 
                           PCBranchD_wire_18_port, PCBranchD(17) => 
                           PCBranchD_wire_17_port, PCBranchD(16) => 
                           PCBranchD_wire_16_port, PCBranchD(15) => 
                           PCBranchD_wire_15_port, PCBranchD(14) => 
                           PCBranchD_wire_14_port, PCBranchD(13) => 
                           PCBranchD_wire_13_port, PCBranchD(12) => 
                           PCBranchD_wire_12_port, PCBranchD(11) => 
                           PCBranchD_wire_11_port, PCBranchD(10) => 
                           PCBranchD_wire_10_port, PCBranchD(9) => 
                           PCBranchD_wire_9_port, PCBranchD(8) => 
                           PCBranchD_wire_8_port, PCBranchD(7) => 
                           PCBranchD_wire_7_port, PCBranchD(6) => 
                           PCBranchD_wire_6_port, PCBranchD(5) => 
                           PCBranchD_wire_5_port, PCBranchD(4) => 
                           PCBranchD_wire_4_port, PCBranchD(3) => 
                           PCBranchD_wire_3_port, PCBranchD(2) => 
                           PCBranchD_wire_2_port, PCBranchD(1) => 
                           PCBranchD_wire_1_port, PCBranchD(0) => 
                           PCBranchD_wire_0_port, PCPlus4F(31) => 
                           PCPlus4F_wire_31_port, PCPlus4F(30) => 
                           PCPlus4F_wire_30_port, PCPlus4F(29) => 
                           PCPlus4F_wire_29_port, PCPlus4F(28) => 
                           PCPlus4F_wire_28_port, PCPlus4F(27) => 
                           PCPlus4F_wire_27_port, PCPlus4F(26) => 
                           PCPlus4F_wire_26_port, PCPlus4F(25) => 
                           PCPlus4F_wire_25_port, PCPlus4F(24) => 
                           PCPlus4F_wire_24_port, PCPlus4F(23) => 
                           PCPlus4F_wire_23_port, PCPlus4F(22) => 
                           PCPlus4F_wire_22_port, PCPlus4F(21) => 
                           PCPlus4F_wire_21_port, PCPlus4F(20) => 
                           PCPlus4F_wire_20_port, PCPlus4F(19) => 
                           PCPlus4F_wire_19_port, PCPlus4F(18) => 
                           PCPlus4F_wire_18_port, PCPlus4F(17) => 
                           PCPlus4F_wire_17_port, PCPlus4F(16) => 
                           PCPlus4F_wire_16_port, PCPlus4F(15) => 
                           PCPlus4F_wire_15_port, PCPlus4F(14) => 
                           PCPlus4F_wire_14_port, PCPlus4F(13) => 
                           PCPlus4F_wire_13_port, PCPlus4F(12) => 
                           PCPlus4F_wire_12_port, PCPlus4F(11) => 
                           PCPlus4F_wire_11_port, PCPlus4F(10) => 
                           PCPlus4F_wire_10_port, PCPlus4F(9) => 
                           PCPlus4F_wire_9_port, PCPlus4F(8) => 
                           PCPlus4F_wire_8_port, PCPlus4F(7) => 
                           PCPlus4F_wire_7_port, PCPlus4F(6) => 
                           PCPlus4F_wire_6_port, PCPlus4F(5) => 
                           PCPlus4F_wire_5_port, PCPlus4F(4) => 
                           PCPlus4F_wire_4_port, PCPlus4F(3) => 
                           PCPlus4F_wire_3_port, PCPlus4F(2) => 
                           PCPlus4F_wire_2_port, PCPlus4F(1) => 
                           PCPlus4F_wire_1_port, PCPlus4F(0) => 
                           PCPlus4F_wire_0_port, InstrD(31) => 
                           InstrD_wire_31_port, InstrD(30) => 
                           InstrD_wire_30_port, InstrD(29) => 
                           InstrD_wire_29_port, InstrD(28) => 
                           InstrD_wire_28_port, InstrD(27) => 
                           InstrD_wire_27_port, InstrD(26) => 
                           InstrD_wire_26_port, InstrD(25) => 
                           InstrD_wire_25_port, InstrD(24) => 
                           InstrD_wire_24_port, InstrD(23) => 
                           InstrD_wire_23_port, InstrD(22) => 
                           InstrD_wire_22_port, InstrD(21) => 
                           InstrD_wire_21_port, InstrD(20) => 
                           InstrD_wire_20_port, InstrD(19) => 
                           InstrD_wire_19_port, InstrD(18) => 
                           InstrD_wire_18_port, InstrD(17) => 
                           InstrD_wire_17_port, InstrD(16) => 
                           InstrD_wire_16_port, InstrD(15) => 
                           InstrD_wire_15_port, InstrD(14) => 
                           InstrD_wire_14_port, InstrD(13) => 
                           InstrD_wire_13_port, InstrD(12) => 
                           InstrD_wire_12_port, InstrD(11) => 
                           InstrD_wire_11_port, InstrD(10) => 
                           InstrD_wire_10_port, InstrD(9) => InstrD_wire_9_port
                           , InstrD(8) => InstrD_wire_8_port, InstrD(7) => 
                           InstrD_wire_7_port, InstrD(6) => InstrD_wire_6_port,
                           InstrD(5) => InstrD_wire_5_port, InstrD(4) => 
                           InstrD_wire_4_port, InstrD(3) => InstrD_wire_3_port,
                           InstrD(2) => InstrD_wire_2_port, InstrD(1) => 
                           InstrD_wire_1_port, InstrD(0) => InstrD_wire_0_port,
                           address_to_iram(31) => address_to_iram(31), 
                           address_to_iram(30) => address_to_iram(30), 
                           address_to_iram(29) => address_to_iram(29), 
                           address_to_iram(28) => address_to_iram(28), 
                           address_to_iram(27) => address_to_iram(27), 
                           address_to_iram(26) => address_to_iram(26), 
                           address_to_iram(25) => address_to_iram(25), 
                           address_to_iram(24) => address_to_iram(24), 
                           address_to_iram(23) => address_to_iram(23), 
                           address_to_iram(22) => address_to_iram(22), 
                           address_to_iram(21) => address_to_iram(21), 
                           address_to_iram(20) => address_to_iram(20), 
                           address_to_iram(19) => address_to_iram(19), 
                           address_to_iram(18) => address_to_iram(18), 
                           address_to_iram(17) => address_to_iram(17), 
                           address_to_iram(16) => address_to_iram(16), 
                           address_to_iram(15) => address_to_iram(15), 
                           address_to_iram(14) => address_to_iram(14), 
                           address_to_iram(13) => address_to_iram(13), 
                           address_to_iram(12) => address_to_iram(12), 
                           address_to_iram(11) => address_to_iram(11), 
                           address_to_iram(10) => address_to_iram(10), 
                           address_to_iram(9) => address_to_iram(9), 
                           address_to_iram(8) => address_to_iram(8), 
                           address_to_iram(7) => address_to_iram(7), 
                           address_to_iram(6) => address_to_iram(6), 
                           address_to_iram(5) => address_to_iram(5), 
                           address_to_iram(4) => address_to_iram(4), 
                           address_to_iram(3) => address_to_iram(3), 
                           address_to_iram(2) => address_to_iram(2), 
                           address_to_iram(1) => address_to_iram(1), 
                           address_to_iram(0) => address_to_iram(0), 
                           iram_to_dlx(31) => iram_to_dlx(31), iram_to_dlx(30) 
                           => iram_to_dlx(30), iram_to_dlx(29) => 
                           iram_to_dlx(29), iram_to_dlx(28) => iram_to_dlx(28),
                           iram_to_dlx(27) => iram_to_dlx(27), iram_to_dlx(26) 
                           => iram_to_dlx(26), iram_to_dlx(25) => 
                           iram_to_dlx(25), iram_to_dlx(24) => iram_to_dlx(24),
                           iram_to_dlx(23) => iram_to_dlx(23), iram_to_dlx(22) 
                           => iram_to_dlx(22), iram_to_dlx(21) => 
                           iram_to_dlx(21), iram_to_dlx(20) => iram_to_dlx(20),
                           iram_to_dlx(19) => iram_to_dlx(19), iram_to_dlx(18) 
                           => iram_to_dlx(18), iram_to_dlx(17) => 
                           iram_to_dlx(17), iram_to_dlx(16) => iram_to_dlx(16),
                           iram_to_dlx(15) => iram_to_dlx(15), iram_to_dlx(14) 
                           => iram_to_dlx(14), iram_to_dlx(13) => 
                           iram_to_dlx(13), iram_to_dlx(12) => iram_to_dlx(12),
                           iram_to_dlx(11) => iram_to_dlx(11), iram_to_dlx(10) 
                           => iram_to_dlx(10), iram_to_dlx(9) => iram_to_dlx(9)
                           , iram_to_dlx(8) => iram_to_dlx(8), iram_to_dlx(7) 
                           => iram_to_dlx(7), iram_to_dlx(6) => iram_to_dlx(6),
                           iram_to_dlx(5) => iram_to_dlx(5), iram_to_dlx(4) => 
                           iram_to_dlx(4), iram_to_dlx(3) => iram_to_dlx(3), 
                           iram_to_dlx(2) => iram_to_dlx(2), iram_to_dlx(1) => 
                           iram_to_dlx(1), iram_to_dlx(0) => iram_to_dlx(0), 
                           PCSrcD => PCSrcD, StallF => StallF, clk => clk, rst 
                           => rst);
   decode_stage : Decode_wrapper port map( instrD(31) => IR_31_port, instrD(30)
                           => IR_30_port, instrD(29) => IR_29_port, instrD(28) 
                           => IR_28_port, instrD(27) => IR_27_port, instrD(26) 
                           => IR_26_port, instrD(25) => IR_25_port, instrD(24) 
                           => IR_24_port, instrD(23) => IR_23_port, instrD(22) 
                           => IR_22_port, instrD(21) => IR_21_port, instrD(20) 
                           => IR_20_port, instrD(19) => IR_19_port, instrD(18) 
                           => IR_18_port, instrD(17) => IR_17_port, instrD(16) 
                           => IR_16_port, instrD(15) => IR_15_port, instrD(14) 
                           => IR_14_port, instrD(13) => IR_13_port, instrD(12) 
                           => IR_12_port, instrD(11) => IR_11_port, instrD(10) 
                           => IR_10_port, instrD(9) => IR_9_port, instrD(8) => 
                           IR_8_port, instrD(7) => IR_7_port, instrD(6) => 
                           IR_6_port, instrD(5) => IR_5_port, instrD(4) => 
                           IR_4_port, instrD(3) => IR_3_port, instrD(2) => 
                           IR_2_port, instrD(1) => IR_1_port, instrD(0) => 
                           IR_0_port, PcPlus4D(31) => PCPlus4_31_port, 
                           PcPlus4D(30) => PCPlus4_30_port, PcPlus4D(29) => 
                           PCPlus4_29_port, PcPlus4D(28) => PCPlus4_28_port, 
                           PcPlus4D(27) => PCPlus4_27_port, PcPlus4D(26) => 
                           PCPlus4_26_port, PcPlus4D(25) => PCPlus4_25_port, 
                           PcPlus4D(24) => PCPlus4_24_port, PcPlus4D(23) => 
                           PCPlus4_23_port, PcPlus4D(22) => PCPlus4_22_port, 
                           PcPlus4D(21) => PCPlus4_21_port, PcPlus4D(20) => 
                           PCPlus4_20_port, PcPlus4D(19) => PCPlus4_19_port, 
                           PcPlus4D(18) => PCPlus4_18_port, PcPlus4D(17) => 
                           PCPlus4_17_port, PcPlus4D(16) => PCPlus4_16_port, 
                           PcPlus4D(15) => PCPlus4_15_port, PcPlus4D(14) => 
                           PCPlus4_14_port, PcPlus4D(13) => PCPlus4_13_port, 
                           PcPlus4D(12) => PCPlus4_12_port, PcPlus4D(11) => 
                           PCPlus4_11_port, PcPlus4D(10) => PCPlus4_10_port, 
                           PcPlus4D(9) => PCPlus4_9_port, PcPlus4D(8) => 
                           PCPlus4_8_port, PcPlus4D(7) => PCPlus4_7_port, 
                           PcPlus4D(6) => PCPlus4_6_port, PcPlus4D(5) => 
                           PCPlus4_5_port, PcPlus4D(4) => PCPlus4_4_port, 
                           PcPlus4D(3) => PCPlus4_3_port, PcPlus4D(2) => 
                           PCPlus4_2_port, PcPlus4D(1) => PCPlus4_1_port, 
                           PcPlus4D(0) => PCPlus4_0_port, select_ext => 
                           Select_ext, ForwardAd => ForwardAD, ForwardBD => 
                           ForwardBD, clk => clk, en => en_RF, rst => rst_RF, 
                           RD1_EN => RD1_EN, RD2_EN => RD2_EN, ALUOutM(31) => 
                           ALUOutMOut_wire_31_port, ALUOutM(30) => 
                           ALUOutMOut_wire_30_port, ALUOutM(29) => 
                           ALUOutMOut_wire_29_port, ALUOutM(28) => 
                           ALUOutMOut_wire_28_port, ALUOutM(27) => 
                           ALUOutMOut_wire_27_port, ALUOutM(26) => 
                           ALUOutMOut_wire_26_port, ALUOutM(25) => 
                           ALUOutMOut_wire_25_port, ALUOutM(24) => 
                           ALUOutMOut_wire_24_port, ALUOutM(23) => 
                           ALUOutMOut_wire_23_port, ALUOutM(22) => 
                           ALUOutMOut_wire_22_port, ALUOutM(21) => 
                           ALUOutMOut_wire_21_port, ALUOutM(20) => 
                           ALUOutMOut_wire_20_port, ALUOutM(19) => 
                           ALUOutMOut_wire_19_port, ALUOutM(18) => 
                           ALUOutMOut_wire_18_port, ALUOutM(17) => 
                           ALUOutMOut_wire_17_port, ALUOutM(16) => 
                           ALUOutMOut_wire_16_port, ALUOutM(15) => 
                           ALUOutMOut_wire_15_port, ALUOutM(14) => 
                           ALUOutMOut_wire_14_port, ALUOutM(13) => 
                           ALUOutMOut_wire_13_port, ALUOutM(12) => 
                           ALUOutMOut_wire_12_port, ALUOutM(11) => 
                           ALUOutMOut_wire_11_port, ALUOutM(10) => 
                           ALUOutMOut_wire_10_port, ALUOutM(9) => 
                           ALUOutMOut_wire_9_port, ALUOutM(8) => 
                           ALUOutMOut_wire_8_port, ALUOutM(7) => 
                           ALUOutMOut_wire_7_port, ALUOutM(6) => 
                           ALUOutMOut_wire_6_port, ALUOutM(5) => 
                           ALUOutMOut_wire_5_port, ALUOutM(4) => 
                           ALUOutMOut_wire_4_port, ALUOutM(3) => 
                           ALUOutMOut_wire_3_port, ALUOutM(2) => 
                           ALUOutMOut_wire_2_port, ALUOutM(1) => 
                           ALUOutMOut_wire_1_port, ALUOutM(0) => 
                           ALUOutMOut_wire_0_port, WriteRegW(4) => 
                           WriteRegWBOut_H_4_port, WriteRegW(3) => 
                           WriteRegWBOut_H_3_port, WriteRegW(2) => 
                           WriteRegWBOut_H_2_port, WriteRegW(1) => 
                           WriteRegWBOut_H_1_port, WriteRegW(0) => 
                           WriteRegWBOut_H_0_port, ResultW(31) => 
                           ResultW_wire_31_port, ResultW(30) => 
                           ResultW_wire_30_port, ResultW(29) => 
                           ResultW_wire_29_port, ResultW(28) => 
                           ResultW_wire_28_port, ResultW(27) => 
                           ResultW_wire_27_port, ResultW(26) => 
                           ResultW_wire_26_port, ResultW(25) => 
                           ResultW_wire_25_port, ResultW(24) => 
                           ResultW_wire_24_port, ResultW(23) => 
                           ResultW_wire_23_port, ResultW(22) => 
                           ResultW_wire_22_port, ResultW(21) => 
                           ResultW_wire_21_port, ResultW(20) => 
                           ResultW_wire_20_port, ResultW(19) => 
                           ResultW_wire_19_port, ResultW(18) => 
                           ResultW_wire_18_port, ResultW(17) => 
                           ResultW_wire_17_port, ResultW(16) => 
                           ResultW_wire_16_port, ResultW(15) => 
                           ResultW_wire_15_port, ResultW(14) => 
                           ResultW_wire_14_port, ResultW(13) => 
                           ResultW_wire_13_port, ResultW(12) => 
                           ResultW_wire_12_port, ResultW(11) => 
                           ResultW_wire_11_port, ResultW(10) => 
                           ResultW_wire_10_port, ResultW(9) => 
                           ResultW_wire_9_port, ResultW(8) => 
                           ResultW_wire_8_port, ResultW(7) => 
                           ResultW_wire_7_port, ResultW(6) => 
                           ResultW_wire_6_port, ResultW(5) => 
                           ResultW_wire_5_port, ResultW(4) => 
                           ResultW_wire_4_port, ResultW(3) => 
                           ResultW_wire_3_port, ResultW(2) => 
                           ResultW_wire_2_port, ResultW(1) => 
                           ResultW_wire_1_port, ResultW(0) => 
                           ResultW_wire_0_port, CALL => CALL, RET => RET, IsJal
                           => isJal, Comp_control(1) => Comp_control(1), 
                           Comp_control(0) => Comp_control(0), RegWriteW => 
                           RegWriteW, Memory_in(31) => X_Logic0_port, 
                           Memory_in(30) => X_Logic0_port, Memory_in(29) => 
                           X_Logic0_port, Memory_in(28) => X_Logic0_port, 
                           Memory_in(27) => X_Logic0_port, Memory_in(26) => 
                           X_Logic0_port, Memory_in(25) => X_Logic0_port, 
                           Memory_in(24) => X_Logic0_port, Memory_in(23) => 
                           X_Logic0_port, Memory_in(22) => X_Logic0_port, 
                           Memory_in(21) => X_Logic0_port, Memory_in(20) => 
                           X_Logic0_port, Memory_in(19) => X_Logic0_port, 
                           Memory_in(18) => X_Logic0_port, Memory_in(17) => 
                           X_Logic0_port, Memory_in(16) => X_Logic0_port, 
                           Memory_in(15) => X_Logic0_port, Memory_in(14) => 
                           X_Logic0_port, Memory_in(13) => X_Logic0_port, 
                           Memory_in(12) => X_Logic0_port, Memory_in(11) => 
                           X_Logic0_port, Memory_in(10) => X_Logic0_port, 
                           Memory_in(9) => X_Logic0_port, Memory_in(8) => 
                           X_Logic0_port, Memory_in(7) => X_Logic0_port, 
                           Memory_in(6) => X_Logic0_port, Memory_in(5) => 
                           X_Logic0_port, Memory_in(4) => X_Logic0_port, 
                           Memory_in(3) => X_Logic0_port, Memory_in(2) => 
                           X_Logic0_port, Memory_in(1) => X_Logic0_port, 
                           Memory_in(0) => X_Logic0_port, Memory_out(31) => 
                           n_1798, Memory_out(30) => n_1799, Memory_out(29) => 
                           n_1800, Memory_out(28) => n_1801, Memory_out(27) => 
                           n_1802, Memory_out(26) => n_1803, Memory_out(25) => 
                           n_1804, Memory_out(24) => n_1805, Memory_out(23) => 
                           n_1806, Memory_out(22) => n_1807, Memory_out(21) => 
                           n_1808, Memory_out(20) => n_1809, Memory_out(19) => 
                           n_1810, Memory_out(18) => n_1811, Memory_out(17) => 
                           n_1812, Memory_out(16) => n_1813, Memory_out(15) => 
                           n_1814, Memory_out(14) => n_1815, Memory_out(13) => 
                           n_1816, Memory_out(12) => n_1817, Memory_out(11) => 
                           n_1818, Memory_out(10) => n_1819, Memory_out(9) => 
                           n_1820, Memory_out(8) => n_1821, Memory_out(7) => 
                           n_1822, Memory_out(6) => n_1823, Memory_out(5) => 
                           n_1824, Memory_out(4) => n_1825, Memory_out(3) => 
                           n_1826, Memory_out(2) => n_1827, Memory_out(1) => 
                           n_1828, Memory_out(0) => n_1829, FILL => FILL, SPILL
                           => n_1830, RsD(4) => RsD_H_4_port, RsD(3) => 
                           RsD_H_3_port, RsD(2) => RsD_H_2_port, RsD(1) => 
                           RsD_H_1_port, RsD(0) => RsD_H_0_port, RtD(4) => 
                           RtD_H_4_port, RtD(3) => RtD_H_3_port, RtD(2) => 
                           RtD_H_2_port, RtD(1) => RtD_H_1_port, RtD(0) => 
                           RtD_H_0_port, RdE(4) => RdD_wire_4_port, RdE(3) => 
                           RdD_wire_3_port, RdE(2) => RdD_wire_2_port, RdE(1) 
                           => RdD_wire_1_port, RdE(0) => RdD_wire_0_port, 
                           SignImmD(31) => SignImmD_wire_31_port, SignImmD(30) 
                           => SignImmD_wire_30_port, SignImmD(29) => 
                           SignImmD_wire_29_port, SignImmD(28) => 
                           SignImmD_wire_28_port, SignImmD(27) => 
                           SignImmD_wire_27_port, SignImmD(26) => 
                           SignImmD_wire_26_port, SignImmD(25) => 
                           SignImmD_wire_25_port, SignImmD(24) => 
                           SignImmD_wire_24_port, SignImmD(23) => 
                           SignImmD_wire_23_port, SignImmD(22) => 
                           SignImmD_wire_22_port, SignImmD(21) => 
                           SignImmD_wire_21_port, SignImmD(20) => 
                           SignImmD_wire_20_port, SignImmD(19) => 
                           SignImmD_wire_19_port, SignImmD(18) => 
                           SignImmD_wire_18_port, SignImmD(17) => 
                           SignImmD_wire_17_port, SignImmD(16) => 
                           SignImmD_wire_16_port, SignImmD(15) => 
                           SignImmD_wire_15_port, SignImmD(14) => 
                           SignImmD_wire_14_port, SignImmD(13) => 
                           SignImmD_wire_13_port, SignImmD(12) => 
                           SignImmD_wire_12_port, SignImmD(11) => 
                           SignImmD_wire_11_port, SignImmD(10) => 
                           SignImmD_wire_10_port, SignImmD(9) => 
                           SignImmD_wire_9_port, SignImmD(8) => 
                           SignImmD_wire_8_port, SignImmD(7) => 
                           SignImmD_wire_7_port, SignImmD(6) => 
                           SignImmD_wire_6_port, SignImmD(5) => 
                           SignImmD_wire_5_port, SignImmD(4) => 
                           SignImmD_wire_4_port, SignImmD(3) => 
                           SignImmD_wire_3_port, SignImmD(2) => 
                           SignImmD_wire_2_port, SignImmD(1) => 
                           SignImmD_wire_1_port, SignImmD(0) => 
                           SignImmD_wire_0_port, PCBranchD(31) => 
                           PCBranchD_wire_31_port, PCBranchD(30) => 
                           PCBranchD_wire_30_port, PCBranchD(29) => 
                           PCBranchD_wire_29_port, PCBranchD(28) => 
                           PCBranchD_wire_28_port, PCBranchD(27) => 
                           PCBranchD_wire_27_port, PCBranchD(26) => 
                           PCBranchD_wire_26_port, PCBranchD(25) => 
                           PCBranchD_wire_25_port, PCBranchD(24) => 
                           PCBranchD_wire_24_port, PCBranchD(23) => 
                           PCBranchD_wire_23_port, PCBranchD(22) => 
                           PCBranchD_wire_22_port, PCBranchD(21) => 
                           PCBranchD_wire_21_port, PCBranchD(20) => 
                           PCBranchD_wire_20_port, PCBranchD(19) => 
                           PCBranchD_wire_19_port, PCBranchD(18) => 
                           PCBranchD_wire_18_port, PCBranchD(17) => 
                           PCBranchD_wire_17_port, PCBranchD(16) => 
                           PCBranchD_wire_16_port, PCBranchD(15) => 
                           PCBranchD_wire_15_port, PCBranchD(14) => 
                           PCBranchD_wire_14_port, PCBranchD(13) => 
                           PCBranchD_wire_13_port, PCBranchD(12) => 
                           PCBranchD_wire_12_port, PCBranchD(11) => 
                           PCBranchD_wire_11_port, PCBranchD(10) => 
                           PCBranchD_wire_10_port, PCBranchD(9) => 
                           PCBranchD_wire_9_port, PCBranchD(8) => 
                           PCBranchD_wire_8_port, PCBranchD(7) => 
                           PCBranchD_wire_7_port, PCBranchD(6) => 
                           PCBranchD_wire_6_port, PCBranchD(5) => 
                           PCBranchD_wire_5_port, PCBranchD(4) => 
                           PCBranchD_wire_4_port, PCBranchD(3) => 
                           PCBranchD_wire_3_port, PCBranchD(2) => 
                           PCBranchD_wire_2_port, PCBranchD(1) => 
                           PCBranchD_wire_1_port, PCBranchD(0) => 
                           PCBranchD_wire_0_port, EqualD => EqualD, OP(5) => 
                           OP(5), OP(4) => OP(4), OP(3) => OP(3), OP(2) => 
                           OP(2), OP(1) => OP(1), OP(0) => OP(0), FUNC(10) => 
                           FUNC(10), FUNC(9) => FUNC(9), FUNC(8) => FUNC(8), 
                           FUNC(7) => FUNC(7), FUNC(6) => FUNC(6), FUNC(5) => 
                           FUNC(5), FUNC(4) => FUNC(4), FUNC(3) => FUNC(3), 
                           FUNC(2) => FUNC(2), FUNC(1) => FUNC(1), FUNC(0) => 
                           FUNC(0), RD1(31) => RD1_wire_31_port, RD1(30) => 
                           RD1_wire_30_port, RD1(29) => RD1_wire_29_port, 
                           RD1(28) => RD1_wire_28_port, RD1(27) => 
                           RD1_wire_27_port, RD1(26) => RD1_wire_26_port, 
                           RD1(25) => RD1_wire_25_port, RD1(24) => 
                           RD1_wire_24_port, RD1(23) => RD1_wire_23_port, 
                           RD1(22) => RD1_wire_22_port, RD1(21) => 
                           RD1_wire_21_port, RD1(20) => RD1_wire_20_port, 
                           RD1(19) => RD1_wire_19_port, RD1(18) => 
                           RD1_wire_18_port, RD1(17) => RD1_wire_17_port, 
                           RD1(16) => RD1_wire_16_port, RD1(15) => 
                           RD1_wire_15_port, RD1(14) => RD1_wire_14_port, 
                           RD1(13) => RD1_wire_13_port, RD1(12) => 
                           RD1_wire_12_port, RD1(11) => RD1_wire_11_port, 
                           RD1(10) => RD1_wire_10_port, RD1(9) => 
                           RD1_wire_9_port, RD1(8) => RD1_wire_8_port, RD1(7) 
                           => RD1_wire_7_port, RD1(6) => RD1_wire_6_port, 
                           RD1(5) => RD1_wire_5_port, RD1(4) => RD1_wire_4_port
                           , RD1(3) => RD1_wire_3_port, RD1(2) => 
                           RD1_wire_2_port, RD1(1) => RD1_wire_1_port, RD1(0) 
                           => RD1_wire_0_port, RD2(31) => RD2_wire_31_port, 
                           RD2(30) => RD2_wire_30_port, RD2(29) => 
                           RD2_wire_29_port, RD2(28) => RD2_wire_28_port, 
                           RD2(27) => RD2_wire_27_port, RD2(26) => 
                           RD2_wire_26_port, RD2(25) => RD2_wire_25_port, 
                           RD2(24) => RD2_wire_24_port, RD2(23) => 
                           RD2_wire_23_port, RD2(22) => RD2_wire_22_port, 
                           RD2(21) => RD2_wire_21_port, RD2(20) => 
                           RD2_wire_20_port, RD2(19) => RD2_wire_19_port, 
                           RD2(18) => RD2_wire_18_port, RD2(17) => 
                           RD2_wire_17_port, RD2(16) => RD2_wire_16_port, 
                           RD2(15) => RD2_wire_15_port, RD2(14) => 
                           RD2_wire_14_port, RD2(13) => RD2_wire_13_port, 
                           RD2(12) => RD2_wire_12_port, RD2(11) => 
                           RD2_wire_11_port, RD2(10) => RD2_wire_10_port, 
                           RD2(9) => RD2_wire_9_port, RD2(8) => RD2_wire_8_port
                           , RD2(7) => RD2_wire_7_port, RD2(6) => 
                           RD2_wire_6_port, RD2(5) => RD2_wire_5_port, RD2(4) 
                           => RD2_wire_4_port, RD2(3) => RD2_wire_3_port, 
                           RD2(2) => RD2_wire_2_port, RD2(1) => RD2_wire_1_port
                           , RD2(0) => RD2_wire_0_port);
   execute_stage : execute_stage_wrapper_NBIT32_N32 port map( en_alu => en_ALU,
                           RD1E(31) => RD1_31_port, RD1E(30) => RD1_30_port, 
                           RD1E(29) => RD1_29_port, RD1E(28) => RD1_28_port, 
                           RD1E(27) => RD1_27_port, RD1E(26) => RD1_26_port, 
                           RD1E(25) => RD1_25_port, RD1E(24) => RD1_24_port, 
                           RD1E(23) => RD1_23_port, RD1E(22) => RD1_22_port, 
                           RD1E(21) => RD1_21_port, RD1E(20) => RD1_20_port, 
                           RD1E(19) => RD1_19_port, RD1E(18) => RD1_18_port, 
                           RD1E(17) => RD1_17_port, RD1E(16) => RD1_16_port, 
                           RD1E(15) => RD1_15_port, RD1E(14) => RD1_14_port, 
                           RD1E(13) => RD1_13_port, RD1E(12) => RD1_12_port, 
                           RD1E(11) => RD1_11_port, RD1E(10) => RD1_10_port, 
                           RD1E(9) => RD1_9_port, RD1E(8) => RD1_8_port, 
                           RD1E(7) => RD1_7_port, RD1E(6) => RD1_6_port, 
                           RD1E(5) => RD1_5_port, RD1E(4) => RD1_4_port, 
                           RD1E(3) => RD1_3_port, RD1E(2) => RD1_2_port, 
                           RD1E(1) => RD1_1_port, RD1E(0) => RD1_0_port, 
                           RD2E(31) => RD2_31_port, RD2E(30) => RD2_30_port, 
                           RD2E(29) => RD2_29_port, RD2E(28) => RD2_28_port, 
                           RD2E(27) => RD2_27_port, RD2E(26) => RD2_26_port, 
                           RD2E(25) => RD2_25_port, RD2E(24) => RD2_24_port, 
                           RD2E(23) => RD2_23_port, RD2E(22) => RD2_22_port, 
                           RD2E(21) => RD2_21_port, RD2E(20) => RD2_20_port, 
                           RD2E(19) => RD2_19_port, RD2E(18) => RD2_18_port, 
                           RD2E(17) => RD2_17_port, RD2E(16) => RD2_16_port, 
                           RD2E(15) => RD2_15_port, RD2E(14) => RD2_14_port, 
                           RD2E(13) => RD2_13_port, RD2E(12) => RD2_12_port, 
                           RD2E(11) => RD2_11_port, RD2E(10) => RD2_10_port, 
                           RD2E(9) => RD2_9_port, RD2E(8) => RD2_8_port, 
                           RD2E(7) => RD2_7_port, RD2E(6) => RD2_6_port, 
                           RD2E(5) => RD2_5_port, RD2E(4) => RD2_4_port, 
                           RD2E(3) => RD2_3_port, RD2E(2) => RD2_2_port, 
                           RD2E(1) => RD2_1_port, RD2E(0) => RD2_0_port, RsE(4)
                           => RsD_4_port, RsE(3) => RsD_3_port, RsE(2) => 
                           RsD_2_port, RsE(1) => RsD_1_port, RsE(0) => 
                           RsD_0_port, RdE(4) => RdD_4_port, RdE(3) => 
                           RdD_3_port, RdE(2) => RdD_2_port, RdE(1) => 
                           RdD_1_port, RdE(0) => RdD_0_port, RtE(4) => 
                           RtD_4_port, RtE(3) => RtD_3_port, RtE(2) => 
                           RtD_2_port, RtE(1) => RtD_1_port, RtE(0) => 
                           RtD_0_port, SignImmE(31) => SignImmD_31_port, 
                           SignImmE(30) => SignImmD_30_port, SignImmE(29) => 
                           SignImmD_29_port, SignImmE(28) => SignImmD_28_port, 
                           SignImmE(27) => SignImmD_27_port, SignImmE(26) => 
                           SignImmD_26_port, SignImmE(25) => SignImmD_25_port, 
                           SignImmE(24) => SignImmD_24_port, SignImmE(23) => 
                           SignImmD_23_port, SignImmE(22) => SignImmD_22_port, 
                           SignImmE(21) => SignImmD_21_port, SignImmE(20) => 
                           SignImmD_20_port, SignImmE(19) => SignImmD_19_port, 
                           SignImmE(18) => SignImmD_18_port, SignImmE(17) => 
                           SignImmD_17_port, SignImmE(16) => SignImmD_16_port, 
                           SignImmE(15) => SignImmD_15_port, SignImmE(14) => 
                           SignImmD_14_port, SignImmE(13) => SignImmD_13_port, 
                           SignImmE(12) => SignImmD_12_port, SignImmE(11) => 
                           SignImmD_11_port, SignImmE(10) => SignImmD_10_port, 
                           SignImmE(9) => SignImmD_9_port, SignImmE(8) => 
                           SignImmD_8_port, SignImmE(7) => SignImmD_7_port, 
                           SignImmE(6) => SignImmD_6_port, SignImmE(5) => 
                           SignImmD_5_port, SignImmE(4) => SignImmD_4_port, 
                           SignImmE(3) => SignImmD_3_port, SignImmE(2) => 
                           SignImmD_2_port, SignImmE(1) => SignImmD_1_port, 
                           SignImmE(0) => SignImmD_0_port, ALUOutME(31) => 
                           ALUOutMOut_wire_31_port, ALUOutME(30) => 
                           ALUOutMOut_wire_30_port, ALUOutME(29) => 
                           ALUOutMOut_wire_29_port, ALUOutME(28) => 
                           ALUOutMOut_wire_28_port, ALUOutME(27) => 
                           ALUOutMOut_wire_27_port, ALUOutME(26) => 
                           ALUOutMOut_wire_26_port, ALUOutME(25) => 
                           ALUOutMOut_wire_25_port, ALUOutME(24) => 
                           ALUOutMOut_wire_24_port, ALUOutME(23) => 
                           ALUOutMOut_wire_23_port, ALUOutME(22) => 
                           ALUOutMOut_wire_22_port, ALUOutME(21) => 
                           ALUOutMOut_wire_21_port, ALUOutME(20) => 
                           ALUOutMOut_wire_20_port, ALUOutME(19) => 
                           ALUOutMOut_wire_19_port, ALUOutME(18) => 
                           ALUOutMOut_wire_18_port, ALUOutME(17) => 
                           ALUOutMOut_wire_17_port, ALUOutME(16) => 
                           ALUOutMOut_wire_16_port, ALUOutME(15) => 
                           ALUOutMOut_wire_15_port, ALUOutME(14) => 
                           ALUOutMOut_wire_14_port, ALUOutME(13) => 
                           ALUOutMOut_wire_13_port, ALUOutME(12) => 
                           ALUOutMOut_wire_12_port, ALUOutME(11) => 
                           ALUOutMOut_wire_11_port, ALUOutME(10) => 
                           ALUOutMOut_wire_10_port, ALUOutME(9) => 
                           ALUOutMOut_wire_9_port, ALUOutME(8) => 
                           ALUOutMOut_wire_8_port, ALUOutME(7) => 
                           ALUOutMOut_wire_7_port, ALUOutME(6) => 
                           ALUOutMOut_wire_6_port, ALUOutME(5) => 
                           ALUOutMOut_wire_5_port, ALUOutME(4) => 
                           ALUOutMOut_wire_4_port, ALUOutME(3) => 
                           ALUOutMOut_wire_3_port, ALUOutME(2) => 
                           ALUOutMOut_wire_2_port, ALUOutME(1) => 
                           ALUOutMOut_wire_1_port, ALUOutME(0) => 
                           ALUOutMOut_wire_0_port, ResultWE(31) => 
                           ResultW_wire_31_port, ResultWE(30) => 
                           ResultW_wire_30_port, ResultWE(29) => 
                           ResultW_wire_29_port, ResultWE(28) => 
                           ResultW_wire_28_port, ResultWE(27) => 
                           ResultW_wire_27_port, ResultWE(26) => 
                           ResultW_wire_26_port, ResultWE(25) => 
                           ResultW_wire_25_port, ResultWE(24) => 
                           ResultW_wire_24_port, ResultWE(23) => 
                           ResultW_wire_23_port, ResultWE(22) => 
                           ResultW_wire_22_port, ResultWE(21) => 
                           ResultW_wire_21_port, ResultWE(20) => 
                           ResultW_wire_20_port, ResultWE(19) => 
                           ResultW_wire_19_port, ResultWE(18) => 
                           ResultW_wire_18_port, ResultWE(17) => 
                           ResultW_wire_17_port, ResultWE(16) => 
                           ResultW_wire_16_port, ResultWE(15) => 
                           ResultW_wire_15_port, ResultWE(14) => 
                           ResultW_wire_14_port, ResultWE(13) => 
                           ResultW_wire_13_port, ResultWE(12) => 
                           ResultW_wire_12_port, ResultWE(11) => 
                           ResultW_wire_11_port, ResultWE(10) => 
                           ResultW_wire_10_port, ResultWE(9) => 
                           ResultW_wire_9_port, ResultWE(8) => 
                           ResultW_wire_8_port, ResultWE(7) => 
                           ResultW_wire_7_port, ResultWE(6) => 
                           ResultW_wire_6_port, ResultWE(5) => 
                           ResultW_wire_5_port, ResultWE(4) => 
                           ResultW_wire_4_port, ResultWE(3) => 
                           ResultW_wire_3_port, ResultWE(2) => 
                           ResultW_wire_2_port, ResultWE(1) => 
                           ResultW_wire_1_port, ResultWE(0) => 
                           ResultW_wire_0_port, ALUoutE(31) => 
                           ALUOutE_wire_31_port, ALUoutE(30) => 
                           ALUOutE_wire_30_port, ALUoutE(29) => 
                           ALUOutE_wire_29_port, ALUoutE(28) => 
                           ALUOutE_wire_28_port, ALUoutE(27) => 
                           ALUOutE_wire_27_port, ALUoutE(26) => 
                           ALUOutE_wire_26_port, ALUoutE(25) => 
                           ALUOutE_wire_25_port, ALUoutE(24) => 
                           ALUOutE_wire_24_port, ALUoutE(23) => 
                           ALUOutE_wire_23_port, ALUoutE(22) => 
                           ALUOutE_wire_22_port, ALUoutE(21) => 
                           ALUOutE_wire_21_port, ALUoutE(20) => 
                           ALUOutE_wire_20_port, ALUoutE(19) => 
                           ALUOutE_wire_19_port, ALUoutE(18) => 
                           ALUOutE_wire_18_port, ALUoutE(17) => 
                           ALUOutE_wire_17_port, ALUoutE(16) => 
                           ALUOutE_wire_16_port, ALUoutE(15) => 
                           ALUOutE_wire_15_port, ALUoutE(14) => 
                           ALUOutE_wire_14_port, ALUoutE(13) => 
                           ALUOutE_wire_13_port, ALUoutE(12) => 
                           ALUOutE_wire_12_port, ALUoutE(11) => 
                           ALUOutE_wire_11_port, ALUoutE(10) => 
                           ALUOutE_wire_10_port, ALUoutE(9) => 
                           ALUOutE_wire_9_port, ALUoutE(8) => 
                           ALUOutE_wire_8_port, ALUoutE(7) => 
                           ALUOutE_wire_7_port, ALUoutE(6) => 
                           ALUOutE_wire_6_port, ALUoutE(5) => 
                           ALUOutE_wire_5_port, ALUoutE(4) => 
                           ALUOutE_wire_4_port, ALUoutE(3) => 
                           ALUOutE_wire_3_port, ALUoutE(2) => 
                           ALUOutE_wire_2_port, ALUoutE(1) => 
                           ALUOutE_wire_1_port, ALUoutE(0) => 
                           ALUOutE_wire_0_port, WriteRegE(4) => 
                           WriteRegE_H_4_port, WriteRegE(3) => 
                           WriteRegE_H_3_port, WriteRegE(2) => 
                           WriteRegE_H_2_port, WriteRegE(1) => 
                           WriteRegE_H_1_port, WriteRegE(0) => 
                           WriteRegE_H_0_port, WriteDataE(31) => 
                           WriteDataE_wire_31_port, WriteDataE(30) => 
                           WriteDataE_wire_30_port, WriteDataE(29) => 
                           WriteDataE_wire_29_port, WriteDataE(28) => 
                           WriteDataE_wire_28_port, WriteDataE(27) => 
                           WriteDataE_wire_27_port, WriteDataE(26) => 
                           WriteDataE_wire_26_port, WriteDataE(25) => 
                           WriteDataE_wire_25_port, WriteDataE(24) => 
                           WriteDataE_wire_24_port, WriteDataE(23) => 
                           WriteDataE_wire_23_port, WriteDataE(22) => 
                           WriteDataE_wire_22_port, WriteDataE(21) => 
                           WriteDataE_wire_21_port, WriteDataE(20) => 
                           WriteDataE_wire_20_port, WriteDataE(19) => 
                           WriteDataE_wire_19_port, WriteDataE(18) => 
                           WriteDataE_wire_18_port, WriteDataE(17) => 
                           WriteDataE_wire_17_port, WriteDataE(16) => 
                           WriteDataE_wire_16_port, WriteDataE(15) => 
                           WriteDataE_wire_15_port, WriteDataE(14) => 
                           WriteDataE_wire_14_port, WriteDataE(13) => 
                           WriteDataE_wire_13_port, WriteDataE(12) => 
                           WriteDataE_wire_12_port, WriteDataE(11) => 
                           WriteDataE_wire_11_port, WriteDataE(10) => 
                           WriteDataE_wire_10_port, WriteDataE(9) => 
                           WriteDataE_wire_9_port, WriteDataE(8) => 
                           WriteDataE_wire_8_port, WriteDataE(7) => 
                           WriteDataE_wire_7_port, WriteDataE(6) => 
                           WriteDataE_wire_6_port, WriteDataE(5) => 
                           WriteDataE_wire_5_port, WriteDataE(4) => 
                           WriteDataE_wire_4_port, WriteDataE(3) => 
                           WriteDataE_wire_3_port, WriteDataE(2) => 
                           WriteDataE_wire_2_port, WriteDataE(1) => 
                           WriteDataE_wire_1_port, WriteDataE(0) => 
                           WriteDataE_wire_0_port, ForwardAE(1) => ForwardAE(1)
                           , ForwardAE(0) => ForwardAE(0), ForwardBE(1) => 
                           ForwardBE(1), ForwardBE(0) => ForwardBE(0), RsE_o(4)
                           => RsE_H(4), RsE_o(3) => RsE_H(3), RsE_o(2) => 
                           RsE_H(2), RsE_o(1) => RsE_H(1), RsE_o(0) => RsE_H(0)
                           , RtE_o(4) => RtE_H(4), RtE_o(3) => RtE_H(3), 
                           RtE_o(2) => RtE_H(2), RtE_o(1) => RtE_H(1), RtE_o(0)
                           => RtE_H(0), RegDstE => RegDstE, ALUSrcE => ALUSrcE,
                           ALUcontrolE(5) => ALUControlE(5), ALUcontrolE(4) => 
                           ALUControlE(4), ALUcontrolE(3) => ALUControlE(3), 
                           ALUcontrolE(2) => ALUControlE(2), ALUcontrolE(1) => 
                           ALUControlE(1), ALUcontrolE(0) => ALUControlE(0));
   memory_stage : memory_unit_nbit32_nwords64 port map( ALUOutMIn(31) => 
                           ALUOutE_31_port, ALUOutMIn(30) => ALUOutE_30_port, 
                           ALUOutMIn(29) => ALUOutE_29_port, ALUOutMIn(28) => 
                           ALUOutE_28_port, ALUOutMIn(27) => ALUOutE_27_port, 
                           ALUOutMIn(26) => ALUOutE_26_port, ALUOutMIn(25) => 
                           ALUOutE_25_port, ALUOutMIn(24) => ALUOutE_24_port, 
                           ALUOutMIn(23) => ALUOutE_23_port, ALUOutMIn(22) => 
                           ALUOutE_22_port, ALUOutMIn(21) => ALUOutE_21_port, 
                           ALUOutMIn(20) => ALUOutE_20_port, ALUOutMIn(19) => 
                           ALUOutE_19_port, ALUOutMIn(18) => ALUOutE_18_port, 
                           ALUOutMIn(17) => ALUOutE_17_port, ALUOutMIn(16) => 
                           ALUOutE_16_port, ALUOutMIn(15) => ALUOutE_15_port, 
                           ALUOutMIn(14) => ALUOutE_14_port, ALUOutMIn(13) => 
                           ALUOutE_13_port, ALUOutMIn(12) => ALUOutE_12_port, 
                           ALUOutMIn(11) => ALUOutE_11_port, ALUOutMIn(10) => 
                           ALUOutE_10_port, ALUOutMIn(9) => ALUOutE_9_port, 
                           ALUOutMIn(8) => ALUOutE_8_port, ALUOutMIn(7) => 
                           ALUOutE_7_port, ALUOutMIn(6) => ALUOutE_6_port, 
                           ALUOutMIn(5) => ALUOutE_5_port, ALUOutMIn(4) => 
                           ALUOutE_4_port, ALUOutMIn(3) => ALUOutE_3_port, 
                           ALUOutMIn(2) => ALUOutE_2_port, ALUOutMIn(1) => 
                           ALUOutE_1_port, ALUOutMIn(0) => ALUOutE_0_port, 
                           WriteDataM(31) => WriteDataE_31_port, WriteDataM(30)
                           => WriteDataE_30_port, WriteDataM(29) => 
                           WriteDataE_29_port, WriteDataM(28) => 
                           WriteDataE_28_port, WriteDataM(27) => 
                           WriteDataE_27_port, WriteDataM(26) => 
                           WriteDataE_26_port, WriteDataM(25) => 
                           WriteDataE_25_port, WriteDataM(24) => 
                           WriteDataE_24_port, WriteDataM(23) => 
                           WriteDataE_23_port, WriteDataM(22) => 
                           WriteDataE_22_port, WriteDataM(21) => 
                           WriteDataE_21_port, WriteDataM(20) => 
                           WriteDataE_20_port, WriteDataM(19) => 
                           WriteDataE_19_port, WriteDataM(18) => 
                           WriteDataE_18_port, WriteDataM(17) => 
                           WriteDataE_17_port, WriteDataM(16) => 
                           WriteDataE_16_port, WriteDataM(15) => 
                           WriteDataE_15_port, WriteDataM(14) => 
                           WriteDataE_14_port, WriteDataM(13) => 
                           WriteDataE_13_port, WriteDataM(12) => 
                           WriteDataE_12_port, WriteDataM(11) => 
                           WriteDataE_11_port, WriteDataM(10) => 
                           WriteDataE_10_port, WriteDataM(9) => 
                           WriteDataE_9_port, WriteDataM(8) => 
                           WriteDataE_8_port, WriteDataM(7) => 
                           WriteDataE_7_port, WriteDataM(6) => 
                           WriteDataE_6_port, WriteDataM(5) => 
                           WriteDataE_5_port, WriteDataM(4) => 
                           WriteDataE_4_port, WriteDataM(3) => 
                           WriteDataE_3_port, WriteDataM(2) => 
                           WriteDataE_2_port, WriteDataM(1) => 
                           WriteDataE_1_port, WriteDataM(0) => 
                           WriteDataE_0_port, ReadDataM(31) => 
                           ReadDataM_wire_31_port, ReadDataM(30) => 
                           ReadDataM_wire_30_port, ReadDataM(29) => 
                           ReadDataM_wire_29_port, ReadDataM(28) => 
                           ReadDataM_wire_28_port, ReadDataM(27) => 
                           ReadDataM_wire_27_port, ReadDataM(26) => 
                           ReadDataM_wire_26_port, ReadDataM(25) => 
                           ReadDataM_wire_25_port, ReadDataM(24) => 
                           ReadDataM_wire_24_port, ReadDataM(23) => 
                           ReadDataM_wire_23_port, ReadDataM(22) => 
                           ReadDataM_wire_22_port, ReadDataM(21) => 
                           ReadDataM_wire_21_port, ReadDataM(20) => 
                           ReadDataM_wire_20_port, ReadDataM(19) => 
                           ReadDataM_wire_19_port, ReadDataM(18) => 
                           ReadDataM_wire_18_port, ReadDataM(17) => 
                           ReadDataM_wire_17_port, ReadDataM(16) => 
                           ReadDataM_wire_16_port, ReadDataM(15) => 
                           ReadDataM_wire_15_port, ReadDataM(14) => 
                           ReadDataM_wire_14_port, ReadDataM(13) => 
                           ReadDataM_wire_13_port, ReadDataM(12) => 
                           ReadDataM_wire_12_port, ReadDataM(11) => 
                           ReadDataM_wire_11_port, ReadDataM(10) => 
                           ReadDataM_wire_10_port, ReadDataM(9) => 
                           ReadDataM_wire_9_port, ReadDataM(8) => 
                           ReadDataM_wire_8_port, ReadDataM(7) => 
                           ReadDataM_wire_7_port, ReadDataM(6) => 
                           ReadDataM_wire_6_port, ReadDataM(5) => 
                           ReadDataM_wire_5_port, ReadDataM(4) => 
                           ReadDataM_wire_4_port, ReadDataM(3) => 
                           ReadDataM_wire_3_port, ReadDataM(2) => 
                           ReadDataM_wire_2_port, ReadDataM(1) => 
                           ReadDataM_wire_1_port, ReadDataM(0) => 
                           ReadDataM_wire_0_port, ALUOutMOut(31) => 
                           ALUOutMOut_wire_31_port, ALUOutMOut(30) => 
                           ALUOutMOut_wire_30_port, ALUOutMOut(29) => 
                           ALUOutMOut_wire_29_port, ALUOutMOut(28) => 
                           ALUOutMOut_wire_28_port, ALUOutMOut(27) => 
                           ALUOutMOut_wire_27_port, ALUOutMOut(26) => 
                           ALUOutMOut_wire_26_port, ALUOutMOut(25) => 
                           ALUOutMOut_wire_25_port, ALUOutMOut(24) => 
                           ALUOutMOut_wire_24_port, ALUOutMOut(23) => 
                           ALUOutMOut_wire_23_port, ALUOutMOut(22) => 
                           ALUOutMOut_wire_22_port, ALUOutMOut(21) => 
                           ALUOutMOut_wire_21_port, ALUOutMOut(20) => 
                           ALUOutMOut_wire_20_port, ALUOutMOut(19) => 
                           ALUOutMOut_wire_19_port, ALUOutMOut(18) => 
                           ALUOutMOut_wire_18_port, ALUOutMOut(17) => 
                           ALUOutMOut_wire_17_port, ALUOutMOut(16) => 
                           ALUOutMOut_wire_16_port, ALUOutMOut(15) => 
                           ALUOutMOut_wire_15_port, ALUOutMOut(14) => 
                           ALUOutMOut_wire_14_port, ALUOutMOut(13) => 
                           ALUOutMOut_wire_13_port, ALUOutMOut(12) => 
                           ALUOutMOut_wire_12_port, ALUOutMOut(11) => 
                           ALUOutMOut_wire_11_port, ALUOutMOut(10) => 
                           ALUOutMOut_wire_10_port, ALUOutMOut(9) => 
                           ALUOutMOut_wire_9_port, ALUOutMOut(8) => 
                           ALUOutMOut_wire_8_port, ALUOutMOut(7) => 
                           ALUOutMOut_wire_7_port, ALUOutMOut(6) => 
                           ALUOutMOut_wire_6_port, ALUOutMOut(5) => 
                           ALUOutMOut_wire_5_port, ALUOutMOut(4) => 
                           ALUOutMOut_wire_4_port, ALUOutMOut(3) => 
                           ALUOutMOut_wire_3_port, ALUOutMOut(2) => 
                           ALUOutMOut_wire_2_port, ALUOutMOut(1) => 
                           ALUOutMOut_wire_1_port, ALUOutMOut(0) => 
                           ALUOutMOut_wire_0_port, address_to_dram(31) => 
                           address_to_dram(31), address_to_dram(30) => 
                           address_to_dram(30), address_to_dram(29) => 
                           address_to_dram(29), address_to_dram(28) => 
                           address_to_dram(28), address_to_dram(27) => 
                           address_to_dram(27), address_to_dram(26) => 
                           address_to_dram(26), address_to_dram(25) => 
                           address_to_dram(25), address_to_dram(24) => 
                           address_to_dram(24), address_to_dram(23) => 
                           address_to_dram(23), address_to_dram(22) => 
                           address_to_dram(22), address_to_dram(21) => 
                           address_to_dram(21), address_to_dram(20) => 
                           address_to_dram(20), address_to_dram(19) => 
                           address_to_dram(19), address_to_dram(18) => 
                           address_to_dram(18), address_to_dram(17) => 
                           address_to_dram(17), address_to_dram(16) => 
                           address_to_dram(16), address_to_dram(15) => 
                           address_to_dram(15), address_to_dram(14) => 
                           address_to_dram(14), address_to_dram(13) => 
                           address_to_dram(13), address_to_dram(12) => 
                           address_to_dram(12), address_to_dram(11) => 
                           address_to_dram(11), address_to_dram(10) => 
                           address_to_dram(10), address_to_dram(9) => 
                           address_to_dram(9), address_to_dram(8) => 
                           address_to_dram(8), address_to_dram(7) => 
                           address_to_dram(7), address_to_dram(6) => 
                           address_to_dram(6), address_to_dram(5) => 
                           address_to_dram(5), address_to_dram(4) => 
                           address_to_dram(4), address_to_dram(3) => 
                           address_to_dram(3), address_to_dram(2) => 
                           address_to_dram(2), address_to_dram(1) => 
                           address_to_dram(1), address_to_dram(0) => 
                           address_to_dram(0), data_to_dram(31) => 
                           data_to_dram(31), data_to_dram(30) => 
                           data_to_dram(30), data_to_dram(29) => 
                           data_to_dram(29), data_to_dram(28) => 
                           data_to_dram(28), data_to_dram(27) => 
                           data_to_dram(27), data_to_dram(26) => 
                           data_to_dram(26), data_to_dram(25) => 
                           data_to_dram(25), data_to_dram(24) => 
                           data_to_dram(24), data_to_dram(23) => 
                           data_to_dram(23), data_to_dram(22) => 
                           data_to_dram(22), data_to_dram(21) => 
                           data_to_dram(21), data_to_dram(20) => 
                           data_to_dram(20), data_to_dram(19) => 
                           data_to_dram(19), data_to_dram(18) => 
                           data_to_dram(18), data_to_dram(17) => 
                           data_to_dram(17), data_to_dram(16) => 
                           data_to_dram(16), data_to_dram(15) => 
                           data_to_dram(15), data_to_dram(14) => 
                           data_to_dram(14), data_to_dram(13) => 
                           data_to_dram(13), data_to_dram(12) => 
                           data_to_dram(12), data_to_dram(11) => 
                           data_to_dram(11), data_to_dram(10) => 
                           data_to_dram(10), data_to_dram(9) => data_to_dram(9)
                           , data_to_dram(8) => data_to_dram(8), 
                           data_to_dram(7) => data_to_dram(7), data_to_dram(6) 
                           => data_to_dram(6), data_to_dram(5) => 
                           data_to_dram(5), data_to_dram(4) => data_to_dram(4),
                           data_to_dram(3) => data_to_dram(3), data_to_dram(2) 
                           => data_to_dram(2), data_to_dram(1) => 
                           data_to_dram(1), data_to_dram(0) => data_to_dram(0),
                           dram_to_dlx(31) => dram_to_dlx(31), dram_to_dlx(30) 
                           => dram_to_dlx(30), dram_to_dlx(29) => 
                           dram_to_dlx(29), dram_to_dlx(28) => dram_to_dlx(28),
                           dram_to_dlx(27) => dram_to_dlx(27), dram_to_dlx(26) 
                           => dram_to_dlx(26), dram_to_dlx(25) => 
                           dram_to_dlx(25), dram_to_dlx(24) => dram_to_dlx(24),
                           dram_to_dlx(23) => dram_to_dlx(23), dram_to_dlx(22) 
                           => dram_to_dlx(22), dram_to_dlx(21) => 
                           dram_to_dlx(21), dram_to_dlx(20) => dram_to_dlx(20),
                           dram_to_dlx(19) => dram_to_dlx(19), dram_to_dlx(18) 
                           => dram_to_dlx(18), dram_to_dlx(17) => 
                           dram_to_dlx(17), dram_to_dlx(16) => dram_to_dlx(16),
                           dram_to_dlx(15) => dram_to_dlx(15), dram_to_dlx(14) 
                           => dram_to_dlx(14), dram_to_dlx(13) => 
                           dram_to_dlx(13), dram_to_dlx(12) => dram_to_dlx(12),
                           dram_to_dlx(11) => dram_to_dlx(11), dram_to_dlx(10) 
                           => dram_to_dlx(10), dram_to_dlx(9) => dram_to_dlx(9)
                           , dram_to_dlx(8) => dram_to_dlx(8), dram_to_dlx(7) 
                           => dram_to_dlx(7), dram_to_dlx(6) => dram_to_dlx(6),
                           dram_to_dlx(5) => dram_to_dlx(5), dram_to_dlx(4) => 
                           dram_to_dlx(4), dram_to_dlx(3) => dram_to_dlx(3), 
                           dram_to_dlx(2) => dram_to_dlx(2), dram_to_dlx(1) => 
                           dram_to_dlx(1), dram_to_dlx(0) => dram_to_dlx(0), 
                           WriteRegMIn(4) => WriteRegE_4_port, WriteRegMIn(3) 
                           => WriteRegE_3_port, WriteRegMIn(2) => 
                           WriteRegE_2_port, WriteRegMIn(1) => WriteRegE_1_port
                           , WriteRegMIn(0) => WriteRegE_0_port, 
                           WriteRegMOut(4) => WriteRegMOut_H_4_port, 
                           WriteRegMOut(3) => WriteRegMOut_H_3_port, 
                           WriteRegMOut(2) => WriteRegMOut_H_2_port, 
                           WriteRegMOut(1) => WriteRegMOut_H_1_port, 
                           WriteRegMOut(0) => WriteRegMOut_H_0_port, clk => clk
                           , rst => rst_mem, MemWriteM => MemWriteM, 
                           MemWriteM_out => dram_we);
   WB_stage : writeback_unit_N32 port map( ReadDataW(31) => ReadDataM_31_port, 
                           ReadDataW(30) => ReadDataM_30_port, ReadDataW(29) =>
                           ReadDataM_29_port, ReadDataW(28) => 
                           ReadDataM_28_port, ReadDataW(27) => 
                           ReadDataM_27_port, ReadDataW(26) => 
                           ReadDataM_26_port, ReadDataW(25) => 
                           ReadDataM_25_port, ReadDataW(24) => 
                           ReadDataM_24_port, ReadDataW(23) => 
                           ReadDataM_23_port, ReadDataW(22) => 
                           ReadDataM_22_port, ReadDataW(21) => 
                           ReadDataM_21_port, ReadDataW(20) => 
                           ReadDataM_20_port, ReadDataW(19) => 
                           ReadDataM_19_port, ReadDataW(18) => 
                           ReadDataM_18_port, ReadDataW(17) => 
                           ReadDataM_17_port, ReadDataW(16) => 
                           ReadDataM_16_port, ReadDataW(15) => 
                           ReadDataM_15_port, ReadDataW(14) => 
                           ReadDataM_14_port, ReadDataW(13) => 
                           ReadDataM_13_port, ReadDataW(12) => 
                           ReadDataM_12_port, ReadDataW(11) => 
                           ReadDataM_11_port, ReadDataW(10) => 
                           ReadDataM_10_port, ReadDataW(9) => ReadDataM_9_port,
                           ReadDataW(8) => ReadDataM_8_port, ReadDataW(7) => 
                           ReadDataM_7_port, ReadDataW(6) => ReadDataM_6_port, 
                           ReadDataW(5) => ReadDataM_5_port, ReadDataW(4) => 
                           ReadDataM_4_port, ReadDataW(3) => ReadDataM_3_port, 
                           ReadDataW(2) => ReadDataM_2_port, ReadDataW(1) => 
                           ReadDataM_1_port, ReadDataW(0) => ReadDataM_0_port, 
                           ALUOutW(31) => ALUOutM_31_port, ALUOutW(30) => 
                           ALUOutM_30_port, ALUOutW(29) => ALUOutM_29_port, 
                           ALUOutW(28) => ALUOutM_28_port, ALUOutW(27) => 
                           ALUOutM_27_port, ALUOutW(26) => ALUOutM_26_port, 
                           ALUOutW(25) => ALUOutM_25_port, ALUOutW(24) => 
                           ALUOutM_24_port, ALUOutW(23) => ALUOutM_23_port, 
                           ALUOutW(22) => ALUOutM_22_port, ALUOutW(21) => 
                           ALUOutM_21_port, ALUOutW(20) => ALUOutM_20_port, 
                           ALUOutW(19) => ALUOutM_19_port, ALUOutW(18) => 
                           ALUOutM_18_port, ALUOutW(17) => ALUOutM_17_port, 
                           ALUOutW(16) => ALUOutM_16_port, ALUOutW(15) => 
                           ALUOutM_15_port, ALUOutW(14) => ALUOutM_14_port, 
                           ALUOutW(13) => ALUOutM_13_port, ALUOutW(12) => 
                           ALUOutM_12_port, ALUOutW(11) => ALUOutM_11_port, 
                           ALUOutW(10) => ALUOutM_10_port, ALUOutW(9) => 
                           ALUOutM_9_port, ALUOutW(8) => ALUOutM_8_port, 
                           ALUOutW(7) => ALUOutM_7_port, ALUOutW(6) => 
                           ALUOutM_6_port, ALUOutW(5) => ALUOutM_5_port, 
                           ALUOutW(4) => ALUOutM_4_port, ALUOutW(3) => 
                           ALUOutM_3_port, ALUOutW(2) => ALUOutM_2_port, 
                           ALUOutW(1) => ALUOutM_1_port, ALUOutW(0) => 
                           ALUOutM_0_port, WriteRegW(4) => WriteRegM_4_port, 
                           WriteRegW(3) => WriteRegM_3_port, WriteRegW(2) => 
                           WriteRegM_2_port, WriteRegW(1) => WriteRegM_1_port, 
                           WriteRegW(0) => WriteRegM_0_port, MemToRegW => 
                           MemToRegW, WriteRegW_out(4) => 
                           WriteRegWBOut_H_4_port, WriteRegW_out(3) => 
                           WriteRegWBOut_H_3_port, WriteRegW_out(2) => 
                           WriteRegWBOut_H_2_port, WriteRegW_out(1) => 
                           WriteRegWBOut_H_1_port, WriteRegW_out(0) => 
                           WriteRegWBOut_H_0_port, ResultW(31) => 
                           ResultW_wire_31_port, ResultW(30) => 
                           ResultW_wire_30_port, ResultW(29) => 
                           ResultW_wire_29_port, ResultW(28) => 
                           ResultW_wire_28_port, ResultW(27) => 
                           ResultW_wire_27_port, ResultW(26) => 
                           ResultW_wire_26_port, ResultW(25) => 
                           ResultW_wire_25_port, ResultW(24) => 
                           ResultW_wire_24_port, ResultW(23) => 
                           ResultW_wire_23_port, ResultW(22) => 
                           ResultW_wire_22_port, ResultW(21) => 
                           ResultW_wire_21_port, ResultW(20) => 
                           ResultW_wire_20_port, ResultW(19) => 
                           ResultW_wire_19_port, ResultW(18) => 
                           ResultW_wire_18_port, ResultW(17) => 
                           ResultW_wire_17_port, ResultW(16) => 
                           ResultW_wire_16_port, ResultW(15) => 
                           ResultW_wire_15_port, ResultW(14) => 
                           ResultW_wire_14_port, ResultW(13) => 
                           ResultW_wire_13_port, ResultW(12) => 
                           ResultW_wire_12_port, ResultW(11) => 
                           ResultW_wire_11_port, ResultW(10) => 
                           ResultW_wire_10_port, ResultW(9) => 
                           ResultW_wire_9_port, ResultW(8) => 
                           ResultW_wire_8_port, ResultW(7) => 
                           ResultW_wire_7_port, ResultW(6) => 
                           ResultW_wire_6_port, ResultW(5) => 
                           ResultW_wire_5_port, ResultW(4) => 
                           ResultW_wire_4_port, ResultW(3) => 
                           ResultW_wire_3_port, ResultW(2) => 
                           ResultW_wire_2_port, ResultW(1) => 
                           ResultW_wire_1_port, ResultW(0) => 
                           ResultW_wire_0_port);
   U3 : OR2_X4 port map( A1 => PCSrcD, A2 => n30, ZN => n28);
   U4 : INV_X4 port map( A => StallD, ZN => n30);
   U5 : CLKBUF_X1 port map( A => n222, Z => n1);
   U6 : CLKBUF_X1 port map( A => n222, Z => n2);
   U7 : CLKBUF_X1 port map( A => n222, Z => n3);
   U8 : CLKBUF_X1 port map( A => n222, Z => n4);
   U9 : CLKBUF_X1 port map( A => n222, Z => n5);
   U10 : CLKBUF_X1 port map( A => n222, Z => n6);
   U11 : CLKBUF_X1 port map( A => n222, Z => n7);
   U12 : CLKBUF_X1 port map( A => n222, Z => n8);
   U13 : CLKBUF_X1 port map( A => n222, Z => n9);
   U14 : CLKBUF_X1 port map( A => n222, Z => n10);
   U15 : CLKBUF_X1 port map( A => n222, Z => n11);
   U16 : CLKBUF_X1 port map( A => n222, Z => n12);
   U17 : CLKBUF_X1 port map( A => n222, Z => n13);
   U18 : CLKBUF_X1 port map( A => n222, Z => n14);
   U19 : CLKBUF_X1 port map( A => n222, Z => n15);
   U20 : CLKBUF_X1 port map( A => n222, Z => n16);
   U21 : CLKBUF_X1 port map( A => n222, Z => n17);
   U22 : CLKBUF_X1 port map( A => n222, Z => n18);
   U23 : CLKBUF_X1 port map( A => n222, Z => n19);
   U24 : CLKBUF_X1 port map( A => n222, Z => n20);
   U25 : CLKBUF_X1 port map( A => n222, Z => n21);
   U26 : CLKBUF_X1 port map( A => n222, Z => n22);
   U27 : CLKBUF_X1 port map( A => n222, Z => n23);
   U28 : CLKBUF_X1 port map( A => n222, Z => n24);
   U29 : CLKBUF_X1 port map( A => n222, Z => n25);
   U30 : CLKBUF_X1 port map( A => n222, Z => n26);
   SPILL <= '0';
   U32 : OAI21_X1 port map( B1 => n94, B2 => n28, A => n29, ZN => n158);
   U33 : NAND2_X1 port map( A1 => PCPlus4F_wire_31_port, A2 => n30, ZN => n29);
   U34 : OAI21_X1 port map( B1 => n95, B2 => n28, A => n31, ZN => n159);
   U35 : NAND2_X1 port map( A1 => PCPlus4F_wire_30_port, A2 => n30, ZN => n31);
   U36 : OAI21_X1 port map( B1 => n96, B2 => n28, A => n32, ZN => n160);
   U37 : NAND2_X1 port map( A1 => PCPlus4F_wire_29_port, A2 => n30, ZN => n32);
   U38 : OAI21_X1 port map( B1 => n97, B2 => n28, A => n33, ZN => n161);
   U39 : NAND2_X1 port map( A1 => PCPlus4F_wire_28_port, A2 => n30, ZN => n33);
   U40 : OAI21_X1 port map( B1 => n98, B2 => n28, A => n34, ZN => n162);
   U41 : NAND2_X1 port map( A1 => PCPlus4F_wire_27_port, A2 => n30, ZN => n34);
   U42 : OAI21_X1 port map( B1 => n99, B2 => n28, A => n35, ZN => n163);
   U43 : NAND2_X1 port map( A1 => PCPlus4F_wire_26_port, A2 => n30, ZN => n35);
   U44 : OAI21_X1 port map( B1 => n100, B2 => n28, A => n36, ZN => n164);
   U45 : NAND2_X1 port map( A1 => PCPlus4F_wire_25_port, A2 => n30, ZN => n36);
   U46 : OAI21_X1 port map( B1 => n101, B2 => n28, A => n37, ZN => n165);
   U47 : NAND2_X1 port map( A1 => PCPlus4F_wire_24_port, A2 => n30, ZN => n37);
   U48 : OAI21_X1 port map( B1 => n102, B2 => n28, A => n38, ZN => n166);
   U49 : NAND2_X1 port map( A1 => PCPlus4F_wire_23_port, A2 => n30, ZN => n38);
   U50 : OAI21_X1 port map( B1 => n103, B2 => n28, A => n39, ZN => n167);
   U51 : NAND2_X1 port map( A1 => PCPlus4F_wire_22_port, A2 => n30, ZN => n39);
   U52 : OAI21_X1 port map( B1 => n104, B2 => n28, A => n40, ZN => n168);
   U53 : NAND2_X1 port map( A1 => PCPlus4F_wire_21_port, A2 => n30, ZN => n40);
   U54 : OAI21_X1 port map( B1 => n105, B2 => n28, A => n41, ZN => n169);
   U55 : NAND2_X1 port map( A1 => PCPlus4F_wire_20_port, A2 => n30, ZN => n41);
   U56 : OAI21_X1 port map( B1 => n106, B2 => n28, A => n42, ZN => n170);
   U57 : NAND2_X1 port map( A1 => PCPlus4F_wire_19_port, A2 => n30, ZN => n42);
   U58 : OAI21_X1 port map( B1 => n107, B2 => n28, A => n43, ZN => n171);
   U59 : NAND2_X1 port map( A1 => PCPlus4F_wire_18_port, A2 => n30, ZN => n43);
   U60 : OAI21_X1 port map( B1 => n108, B2 => n28, A => n44, ZN => n172);
   U61 : NAND2_X1 port map( A1 => PCPlus4F_wire_17_port, A2 => n30, ZN => n44);
   U62 : OAI21_X1 port map( B1 => n109, B2 => n28, A => n45, ZN => n173);
   U63 : NAND2_X1 port map( A1 => PCPlus4F_wire_16_port, A2 => n30, ZN => n45);
   U64 : OAI21_X1 port map( B1 => n110, B2 => n28, A => n46, ZN => n174);
   U65 : NAND2_X1 port map( A1 => PCPlus4F_wire_15_port, A2 => n30, ZN => n46);
   U66 : OAI21_X1 port map( B1 => n111, B2 => n28, A => n47, ZN => n175);
   U67 : NAND2_X1 port map( A1 => PCPlus4F_wire_14_port, A2 => n30, ZN => n47);
   U68 : OAI21_X1 port map( B1 => n112, B2 => n28, A => n48, ZN => n176);
   U69 : NAND2_X1 port map( A1 => PCPlus4F_wire_13_port, A2 => n30, ZN => n48);
   U70 : OAI21_X1 port map( B1 => n113, B2 => n28, A => n49, ZN => n177);
   U71 : NAND2_X1 port map( A1 => PCPlus4F_wire_12_port, A2 => n30, ZN => n49);
   U72 : OAI21_X1 port map( B1 => n114, B2 => n28, A => n50, ZN => n178);
   U73 : NAND2_X1 port map( A1 => PCPlus4F_wire_11_port, A2 => n30, ZN => n50);
   U74 : OAI21_X1 port map( B1 => n115, B2 => n28, A => n51, ZN => n179);
   U75 : NAND2_X1 port map( A1 => PCPlus4F_wire_10_port, A2 => n30, ZN => n51);
   U76 : OAI21_X1 port map( B1 => n116, B2 => n28, A => n52, ZN => n180);
   U77 : NAND2_X1 port map( A1 => PCPlus4F_wire_9_port, A2 => n30, ZN => n52);
   U78 : OAI21_X1 port map( B1 => n117, B2 => n28, A => n53, ZN => n181);
   U79 : NAND2_X1 port map( A1 => PCPlus4F_wire_8_port, A2 => n30, ZN => n53);
   U80 : OAI21_X1 port map( B1 => n118, B2 => n28, A => n54, ZN => n182);
   U81 : NAND2_X1 port map( A1 => PCPlus4F_wire_7_port, A2 => n30, ZN => n54);
   U82 : OAI21_X1 port map( B1 => n119, B2 => n28, A => n55, ZN => n183);
   U83 : NAND2_X1 port map( A1 => PCPlus4F_wire_6_port, A2 => n30, ZN => n55);
   U84 : OAI21_X1 port map( B1 => n120, B2 => n28, A => n56, ZN => n184);
   U85 : NAND2_X1 port map( A1 => PCPlus4F_wire_5_port, A2 => n30, ZN => n56);
   U86 : OAI21_X1 port map( B1 => n121, B2 => n28, A => n57, ZN => n185);
   U87 : NAND2_X1 port map( A1 => PCPlus4F_wire_4_port, A2 => n30, ZN => n57);
   U88 : OAI21_X1 port map( B1 => n122, B2 => n28, A => n58, ZN => n186);
   U89 : NAND2_X1 port map( A1 => PCPlus4F_wire_3_port, A2 => n30, ZN => n58);
   U90 : OAI21_X1 port map( B1 => n123, B2 => n28, A => n59, ZN => n187);
   U91 : NAND2_X1 port map( A1 => PCPlus4F_wire_2_port, A2 => n30, ZN => n59);
   U92 : OAI21_X1 port map( B1 => n124, B2 => n28, A => n60, ZN => n188);
   U93 : NAND2_X1 port map( A1 => PCPlus4F_wire_1_port, A2 => n30, ZN => n60);
   U94 : OAI21_X1 port map( B1 => n125, B2 => n28, A => n61, ZN => n189);
   U95 : NAND2_X1 port map( A1 => PCPlus4F_wire_0_port, A2 => n30, ZN => n61);
   U96 : OAI21_X1 port map( B1 => n157, B2 => n28, A => n62, ZN => n190);
   U97 : NAND2_X1 port map( A1 => InstrD_wire_0_port, A2 => n30, ZN => n62);
   U98 : OAI21_X1 port map( B1 => n156, B2 => n28, A => n63, ZN => n191);
   U99 : NAND2_X1 port map( A1 => InstrD_wire_1_port, A2 => n30, ZN => n63);
   U100 : OAI21_X1 port map( B1 => n155, B2 => n28, A => n64, ZN => n192);
   U101 : NAND2_X1 port map( A1 => InstrD_wire_2_port, A2 => n30, ZN => n64);
   U102 : OAI21_X1 port map( B1 => n154, B2 => n28, A => n65, ZN => n193);
   U103 : NAND2_X1 port map( A1 => InstrD_wire_3_port, A2 => n30, ZN => n65);
   U104 : OAI21_X1 port map( B1 => n153, B2 => n28, A => n66, ZN => n194);
   U105 : NAND2_X1 port map( A1 => InstrD_wire_4_port, A2 => n30, ZN => n66);
   U106 : OAI21_X1 port map( B1 => n152, B2 => n28, A => n67, ZN => n195);
   U107 : NAND2_X1 port map( A1 => InstrD_wire_5_port, A2 => n30, ZN => n67);
   U108 : OAI21_X1 port map( B1 => n151, B2 => n28, A => n68, ZN => n196);
   U109 : NAND2_X1 port map( A1 => InstrD_wire_6_port, A2 => n30, ZN => n68);
   U110 : OAI21_X1 port map( B1 => n150, B2 => n28, A => n69, ZN => n197);
   U111 : NAND2_X1 port map( A1 => InstrD_wire_7_port, A2 => n30, ZN => n69);
   U112 : OAI21_X1 port map( B1 => n149, B2 => n28, A => n70, ZN => n198);
   U113 : NAND2_X1 port map( A1 => InstrD_wire_8_port, A2 => n30, ZN => n70);
   U114 : OAI21_X1 port map( B1 => n148, B2 => n28, A => n71, ZN => n199);
   U115 : NAND2_X1 port map( A1 => InstrD_wire_9_port, A2 => n30, ZN => n71);
   U116 : OAI21_X1 port map( B1 => n147, B2 => n28, A => n72, ZN => n200);
   U117 : NAND2_X1 port map( A1 => InstrD_wire_10_port, A2 => n30, ZN => n72);
   U118 : OAI21_X1 port map( B1 => n146, B2 => n28, A => n73, ZN => n201);
   U119 : NAND2_X1 port map( A1 => InstrD_wire_11_port, A2 => n30, ZN => n73);
   U120 : OAI21_X1 port map( B1 => n145, B2 => n28, A => n74, ZN => n202);
   U121 : NAND2_X1 port map( A1 => InstrD_wire_12_port, A2 => n30, ZN => n74);
   U122 : OAI21_X1 port map( B1 => n144, B2 => n28, A => n75, ZN => n203);
   U123 : NAND2_X1 port map( A1 => InstrD_wire_13_port, A2 => n30, ZN => n75);
   U124 : OAI21_X1 port map( B1 => n143, B2 => n28, A => n76, ZN => n204);
   U125 : NAND2_X1 port map( A1 => InstrD_wire_14_port, A2 => n30, ZN => n76);
   U126 : OAI21_X1 port map( B1 => n142, B2 => n28, A => n77, ZN => n205);
   U127 : NAND2_X1 port map( A1 => InstrD_wire_15_port, A2 => n30, ZN => n77);
   U128 : OAI21_X1 port map( B1 => n141, B2 => n28, A => n78, ZN => n206);
   U129 : NAND2_X1 port map( A1 => InstrD_wire_16_port, A2 => n30, ZN => n78);
   U130 : OAI21_X1 port map( B1 => n140, B2 => n28, A => n79, ZN => n207);
   U131 : NAND2_X1 port map( A1 => InstrD_wire_17_port, A2 => n30, ZN => n79);
   U132 : OAI21_X1 port map( B1 => n139, B2 => n28, A => n80, ZN => n208);
   U133 : NAND2_X1 port map( A1 => InstrD_wire_18_port, A2 => n30, ZN => n80);
   U134 : OAI21_X1 port map( B1 => n138, B2 => n28, A => n81, ZN => n209);
   U135 : NAND2_X1 port map( A1 => InstrD_wire_19_port, A2 => n30, ZN => n81);
   U136 : OAI21_X1 port map( B1 => n137, B2 => n28, A => n82, ZN => n210);
   U137 : NAND2_X1 port map( A1 => InstrD_wire_20_port, A2 => n30, ZN => n82);
   U138 : OAI21_X1 port map( B1 => n136, B2 => n28, A => n83, ZN => n211);
   U139 : NAND2_X1 port map( A1 => InstrD_wire_21_port, A2 => n30, ZN => n83);
   U140 : OAI21_X1 port map( B1 => n135, B2 => n28, A => n84, ZN => n212);
   U141 : NAND2_X1 port map( A1 => InstrD_wire_22_port, A2 => n30, ZN => n84);
   U142 : OAI21_X1 port map( B1 => n134, B2 => n28, A => n85, ZN => n213);
   U143 : NAND2_X1 port map( A1 => InstrD_wire_23_port, A2 => n30, ZN => n85);
   U144 : OAI21_X1 port map( B1 => n133, B2 => n28, A => n86, ZN => n214);
   U145 : NAND2_X1 port map( A1 => InstrD_wire_24_port, A2 => n30, ZN => n86);
   U146 : OAI21_X1 port map( B1 => n132, B2 => n28, A => n87, ZN => n215);
   U147 : NAND2_X1 port map( A1 => InstrD_wire_25_port, A2 => n30, ZN => n87);
   U148 : OAI21_X1 port map( B1 => n131, B2 => n28, A => n88, ZN => n216);
   U149 : NAND2_X1 port map( A1 => InstrD_wire_26_port, A2 => n30, ZN => n88);
   U150 : OAI21_X1 port map( B1 => n130, B2 => n28, A => n89, ZN => n217);
   U151 : NAND2_X1 port map( A1 => InstrD_wire_27_port, A2 => n30, ZN => n89);
   U152 : OAI21_X1 port map( B1 => n129, B2 => n28, A => n90, ZN => n218);
   U153 : NAND2_X1 port map( A1 => InstrD_wire_28_port, A2 => n30, ZN => n90);
   U154 : OAI21_X1 port map( B1 => n128, B2 => n28, A => n91, ZN => n219);
   U155 : NAND2_X1 port map( A1 => InstrD_wire_29_port, A2 => n30, ZN => n91);
   U156 : OAI21_X1 port map( B1 => n127, B2 => n28, A => n92, ZN => n220);
   U157 : NAND2_X1 port map( A1 => InstrD_wire_30_port, A2 => n30, ZN => n92);
   U158 : OAI21_X1 port map( B1 => n126, B2 => n28, A => n93, ZN => n221);
   U159 : NAND2_X1 port map( A1 => InstrD_wire_31_port, A2 => n30, ZN => n93);
   U160 : INV_X1 port map( A => rst, ZN => n222);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity CU_wrapper is

   port( clock, reset : in std_logic;  OPCODE : in std_logic_vector (5 downto 
         0);  FUNC : in std_logic_vector (10 downto 0);  EqualD, FlushE : in 
         std_logic;  PC_SrcD, Select_ext, IsJal, RD1, RD2 : out std_logic;  
         Comp_control : out std_logic_vector (1 downto 0);  ALUcontrolE : out 
         std_logic_vector (5 downto 0);  RegDestE, ALUSrcE, en_ALU, MemWriteM, 
         RegWriteW, MemToRegW, BranchD_H, MemToRegE_H, RegWriteE_H, MemToRegM_H
         , RegWriteM_H, RegWriteW_H, CALL, RET : out std_logic;  FILL, SPILL : 
         in std_logic);

end CU_wrapper;

architecture SYN_Behavioral of CU_wrapper is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component cu
      port( Rst : in std_logic;  OPCODE : in std_logic_vector (5 downto 0);  
            FUNC : in std_logic_vector (10 downto 0);  BranchD, Select_ext, 
            IsJal, RD1, RD2, RegWriteD : out std_logic;  Comp_control : out 
            std_logic_vector (1 downto 0);  en_ALU, RegDestD, ALUSrcD : out 
            std_logic;  ALUcontrolD : out std_logic_vector (5 downto 0);  
            MemWriteD, MemToRegD, CALL, RET : out std_logic;  FILL, SPILL : in 
            std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal MemWriteM_port, RegWriteW_port, MemToRegW_port, MemToRegE_H_port, 
      RegWriteE_H_port, RegWriteM_H_port, n12, n13, n14, n15, n16, n1, n2, n4, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857 : 
      std_logic;

begin
   MemWriteM <= MemWriteM_port;
   RegWriteW <= RegWriteW_port;
   MemToRegW <= MemToRegW_port;
   MemToRegE_H <= MemToRegE_H_port;
   RegWriteE_H <= RegWriteE_H_port;
   MemToRegM_H <= MemWriteM_port;
   RegWriteM_H <= RegWriteM_H_port;
   RegWriteW_H <= RegWriteW_port;
   
   RegWriteE_reg_reg : DFFR_X1 port map( D => n16, CK => clock, RN => n4, Q => 
                           RegWriteM_H_port, QN => n_1832);
   MemWriteE_reg_reg : DFFR_X1 port map( D => n15, CK => clock, RN => n4, Q => 
                           MemWriteM_port, QN => n_1833);
   MemToRegE_reg_reg : DFFR_X1 port map( D => n14, CK => clock, RN => n4, Q => 
                           n1, QN => n_1834);
   RegWriteM_reg_reg : DFFR_X1 port map( D => n12, CK => clock, RN => n4, Q => 
                           RegWriteW_port, QN => n_1835);
   Control : cu port map( Rst => reset, OPCODE(5) => OPCODE(5), OPCODE(4) => 
                           OPCODE(4), OPCODE(3) => OPCODE(3), OPCODE(2) => 
                           OPCODE(2), OPCODE(1) => OPCODE(1), OPCODE(0) => 
                           OPCODE(0), FUNC(10) => FUNC(10), FUNC(9) => FUNC(9),
                           FUNC(8) => FUNC(8), FUNC(7) => FUNC(7), FUNC(6) => 
                           FUNC(6), FUNC(5) => FUNC(5), FUNC(4) => FUNC(4), 
                           FUNC(3) => FUNC(3), FUNC(2) => FUNC(2), FUNC(1) => 
                           FUNC(1), FUNC(0) => FUNC(0), BranchD => n_1836, 
                           Select_ext => n_1837, IsJal => n_1838, RD1 => n_1839
                           , RD2 => n_1840, RegWriteD => n_1841, 
                           Comp_control(1) => n_1842, Comp_control(0) => n_1843
                           , en_ALU => n_1844, RegDestD => n_1845, ALUSrcD => 
                           n_1846, ALUcontrolD(5) => n_1847, ALUcontrolD(4) => 
                           n_1848, ALUcontrolD(3) => n_1849, ALUcontrolD(2) => 
                           n_1850, ALUcontrolD(1) => n_1851, ALUcontrolD(0) => 
                           n_1852, MemWriteD => n_1853, MemToRegD => n_1854, 
                           CALL => n_1855, RET => n_1856, FILL => FILL, SPILL 
                           => SPILL);
   MemToRegM_reg_reg : DFFR_X2 port map( D => n13, CK => clock, RN => n4, Q => 
                           MemToRegW_port, QN => n_1857);
   U3 : MUX2_X1 port map( A => MemToRegE_H_port, B => n1, S => FlushE, Z => n14
                           );
   U4 : MUX2_X1 port map( A => n2, B => MemWriteM_port, S => FlushE, Z => n15);
   U5 : MUX2_X1 port map( A => RegWriteE_H_port, B => RegWriteM_H_port, S => 
                           FlushE, Z => n16);
   RegWriteE_H_port <= '0';
   RegDestE <= '0';
   ALUSrcE <= '0';
   ALUcontrolE(5) <= '0';
   ALUcontrolE(4) <= '0';
   ALUcontrolE(3) <= '0';
   ALUcontrolE(2) <= '0';
   ALUcontrolE(1) <= '0';
   ALUcontrolE(0) <= '0';
   n2 <= '0';
   MemToRegE_H_port <= '0';
   en_ALU <= '0';
   U18 : INV_X1 port map( A => reset, ZN => n4);
   U19 : MUX2_X1 port map( A => n1, B => MemToRegW_port, S => FlushE, Z => n13)
                           ;
   U20 : MUX2_X1 port map( A => RegWriteM_H_port, B => RegWriteW_port, S => 
                           FlushE, Z => n12);
   PC_SrcD <= '0';
   RET <= '0';
   CALL <= '0';
   Comp_control(0) <= '0';
   Comp_control(1) <= '0';
   RD2 <= '0';
   RD1 <= '0';
   IsJal <= '0';
   Select_ext <= '0';
   BranchD_H <= '0';

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nwords64_isize32.all;

entity DLX_nwords64_isize32 is

   port( clk, rst : in std_logic);

end DLX_nwords64_isize32;

architecture SYN_Behavioral of DLX_nwords64_isize32 is

   component hazard_detection_unit
      port( RsD, RtD, RsE, RtE, WriteRegM, WriteRegW, WriteRegE : in 
            std_logic_vector (4 downto 0);  BranchD, MemToRegE, MemToRegM, 
            RegWriteM, RegWriteW, RegWriteE : in std_logic;  ForwardAD, 
            ForwardBD : out std_logic;  ForwardAE, ForwardBE : out 
            std_logic_vector (1 downto 0);  StallF, StallD, FlushE : out 
            std_logic);
   end component;
   
   component DataPath_wrapper
      port( clk, rst : in std_logic;  address_to_iram : out std_logic_vector 
            (31 downto 0);  iram_to_dlx : in std_logic_vector (31 downto 0);  
            address_to_dram, data_to_dram : out std_logic_vector (31 downto 0);
            dram_to_dlx : in std_logic_vector (31 downto 0);  dram_we : out 
            std_logic;  StallF, StallD, ForwardAD, ForwardBD, FlushE, rst_RF, 
            en_RF : in std_logic;  RsD_H, RtD_H : out std_logic_vector (4 
            downto 0);  ForwardAE, ForwardBE : in std_logic_vector (1 downto 0)
            ;  WriteRegE_H, RsE_H, RtE_H, WriteRegMOut_H : out std_logic_vector
            (4 downto 0);  rst_mem : in std_logic;  WriteRegWBOut_H : out 
            std_logic_vector (4 downto 0);  OP : out std_logic_vector (5 downto
            0);  FUNC : out std_logic_vector (10 downto 0);  EqualD, FILL, 
            SPILL : out std_logic;  PCSrcD, RegWriteW, Select_ext, CALL, RET, 
            RD1_EN, RD2_EN, isJal : in std_logic;  Comp_control : in 
            std_logic_vector (1 downto 0);  RegDstE, ALUSrcE : in std_logic;  
            ALUControlE : in std_logic_vector (5 downto 0);  en_ALU, MemWriteM,
            MemToRegW : in std_logic);
   end component;
   
   component CU_wrapper
      port( clock, reset : in std_logic;  OPCODE : in std_logic_vector (5 
            downto 0);  FUNC : in std_logic_vector (10 downto 0);  EqualD, 
            FlushE : in std_logic;  PC_SrcD, Select_ext, IsJal, RD1, RD2 : out 
            std_logic;  Comp_control : out std_logic_vector (1 downto 0);  
            ALUcontrolE : out std_logic_vector (5 downto 0);  RegDestE, ALUSrcE
            , en_ALU, MemWriteM, RegWriteW, MemToRegW, BranchD_H, MemToRegE_H, 
            RegWriteE_H, MemToRegM_H, RegWriteM_H, RegWriteW_H, CALL, RET : out
            std_logic;  FILL, SPILL : in std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, OP_DP_5_port, OP_DP_4_port, 
      OP_DP_3_port, OP_DP_2_port, OP_DP_1_port, OP_DP_0_port, FUNC_DP_10_port, 
      FUNC_DP_9_port, FUNC_DP_8_port, FUNC_DP_7_port, FUNC_DP_6_port, 
      FUNC_DP_5_port, FUNC_DP_4_port, FUNC_DP_3_port, FUNC_DP_2_port, 
      FUNC_DP_1_port, FUNC_DP_0_port, EqualD_DP, FlushE_DP, MemWriteM_CU, 
      RegWriteW_CU, MemToRegW_CU, MemToRegM_H_CU, RegWriteM_H_CU, 
      RegWriteW_H_CU, StallF_DP, StallD_DP, ForwardAD_DP, ForwardBD_DP, 
      RsD_H_DP_4_port, RsD_H_DP_3_port, RsD_H_DP_2_port, RsD_H_DP_1_port, 
      RsD_H_DP_0_port, RtD_H_DP_4_port, RtD_H_DP_3_port, RtD_H_DP_2_port, 
      RtD_H_DP_1_port, RtD_H_DP_0_port, ForwardAE_DP_1_port, 
      ForwardAE_DP_0_port, ForwardBE_DP_1_port, ForwardBE_DP_0_port, 
      WriteRegE_H_DP_4_port, WriteRegE_H_DP_3_port, WriteRegE_H_DP_2_port, 
      WriteRegE_H_DP_1_port, WriteRegE_H_DP_0_port, RsE_H_DP_4_port, 
      RsE_H_DP_3_port, RsE_H_DP_2_port, RsE_H_DP_1_port, RsE_H_DP_0_port, 
      RtE_H_DP_4_port, RtE_H_DP_3_port, RtE_H_DP_2_port, RtE_H_DP_1_port, 
      RtE_H_DP_0_port, WriteRegMOut_H_DP_4_port, WriteRegMOut_H_DP_3_port, 
      WriteRegMOut_H_DP_2_port, WriteRegMOut_H_DP_1_port, 
      WriteRegMOut_H_DP_0_port, WriteRegWBOut_H_DP_4_port, 
      WriteRegWBOut_H_DP_3_port, WriteRegWBOut_H_DP_2_port, 
      WriteRegWBOut_H_DP_1_port, WriteRegWBOut_H_DP_0_port, n1, n2, n_1000, 
      n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   Control_unit : CU_wrapper port map( clock => clk, reset => rst, OPCODE(5) =>
                           OP_DP_5_port, OPCODE(4) => OP_DP_4_port, OPCODE(3) 
                           => OP_DP_3_port, OPCODE(2) => OP_DP_2_port, 
                           OPCODE(1) => OP_DP_1_port, OPCODE(0) => OP_DP_0_port
                           , FUNC(10) => FUNC_DP_10_port, FUNC(9) => 
                           FUNC_DP_9_port, FUNC(8) => FUNC_DP_8_port, FUNC(7) 
                           => FUNC_DP_7_port, FUNC(6) => FUNC_DP_6_port, 
                           FUNC(5) => FUNC_DP_5_port, FUNC(4) => FUNC_DP_4_port
                           , FUNC(3) => FUNC_DP_3_port, FUNC(2) => 
                           FUNC_DP_2_port, FUNC(1) => FUNC_DP_1_port, FUNC(0) 
                           => FUNC_DP_0_port, EqualD => EqualD_DP, FlushE => 
                           FlushE_DP, PC_SrcD => n_1000, Select_ext => n_1001, 
                           IsJal => n_1002, RD1 => n_1003, RD2 => n_1004, 
                           Comp_control(1) => n_1005, Comp_control(0) => n_1006
                           , ALUcontrolE(5) => n_1007, ALUcontrolE(4) => n_1008
                           , ALUcontrolE(3) => n_1009, ALUcontrolE(2) => n_1010
                           , ALUcontrolE(1) => n_1011, ALUcontrolE(0) => n_1012
                           , RegDestE => n_1013, ALUSrcE => n_1014, en_ALU => 
                           n_1015, MemWriteM => MemWriteM_CU, RegWriteW => 
                           RegWriteW_CU, MemToRegW => MemToRegW_CU, BranchD_H 
                           => n_1016, MemToRegE_H => n_1017, RegWriteE_H => 
                           n_1018, MemToRegM_H => MemToRegM_H_CU, RegWriteM_H 
                           => RegWriteM_H_CU, RegWriteW_H => RegWriteW_H_CU, 
                           CALL => n_1019, RET => n_1020, FILL => X_Logic0_port
                           , SPILL => X_Logic0_port);
   DataPath : DataPath_wrapper port map( clk => clk, rst => rst, 
                           address_to_iram(31) => n_1021, address_to_iram(30) 
                           => n_1022, address_to_iram(29) => n_1023, 
                           address_to_iram(28) => n_1024, address_to_iram(27) 
                           => n_1025, address_to_iram(26) => n_1026, 
                           address_to_iram(25) => n_1027, address_to_iram(24) 
                           => n_1028, address_to_iram(23) => n_1029, 
                           address_to_iram(22) => n_1030, address_to_iram(21) 
                           => n_1031, address_to_iram(20) => n_1032, 
                           address_to_iram(19) => n_1033, address_to_iram(18) 
                           => n_1034, address_to_iram(17) => n_1035, 
                           address_to_iram(16) => n_1036, address_to_iram(15) 
                           => n_1037, address_to_iram(14) => n_1038, 
                           address_to_iram(13) => n_1039, address_to_iram(12) 
                           => n_1040, address_to_iram(11) => n_1041, 
                           address_to_iram(10) => n_1042, address_to_iram(9) =>
                           n_1043, address_to_iram(8) => n_1044, 
                           address_to_iram(7) => n_1045, address_to_iram(6) => 
                           n_1046, address_to_iram(5) => n_1047, 
                           address_to_iram(4) => n_1048, address_to_iram(3) => 
                           n_1049, address_to_iram(2) => n_1050, 
                           address_to_iram(1) => n_1051, address_to_iram(0) => 
                           n_1052, iram_to_dlx(31) => X_Logic0_port, 
                           iram_to_dlx(30) => X_Logic0_port, iram_to_dlx(29) =>
                           X_Logic0_port, iram_to_dlx(28) => X_Logic0_port, 
                           iram_to_dlx(27) => X_Logic0_port, iram_to_dlx(26) =>
                           X_Logic0_port, iram_to_dlx(25) => X_Logic0_port, 
                           iram_to_dlx(24) => X_Logic0_port, iram_to_dlx(23) =>
                           X_Logic0_port, iram_to_dlx(22) => X_Logic0_port, 
                           iram_to_dlx(21) => X_Logic0_port, iram_to_dlx(20) =>
                           X_Logic0_port, iram_to_dlx(19) => X_Logic0_port, 
                           iram_to_dlx(18) => X_Logic0_port, iram_to_dlx(17) =>
                           X_Logic0_port, iram_to_dlx(16) => X_Logic0_port, 
                           iram_to_dlx(15) => X_Logic0_port, iram_to_dlx(14) =>
                           X_Logic0_port, iram_to_dlx(13) => X_Logic0_port, 
                           iram_to_dlx(12) => X_Logic0_port, iram_to_dlx(11) =>
                           X_Logic0_port, iram_to_dlx(10) => X_Logic0_port, 
                           iram_to_dlx(9) => X_Logic0_port, iram_to_dlx(8) => 
                           X_Logic0_port, iram_to_dlx(7) => X_Logic0_port, 
                           iram_to_dlx(6) => X_Logic0_port, iram_to_dlx(5) => 
                           X_Logic0_port, iram_to_dlx(4) => X_Logic0_port, 
                           iram_to_dlx(3) => X_Logic0_port, iram_to_dlx(2) => 
                           X_Logic0_port, iram_to_dlx(1) => X_Logic0_port, 
                           iram_to_dlx(0) => X_Logic0_port, address_to_dram(31)
                           => n_1053, address_to_dram(30) => n_1054, 
                           address_to_dram(29) => n_1055, address_to_dram(28) 
                           => n_1056, address_to_dram(27) => n_1057, 
                           address_to_dram(26) => n_1058, address_to_dram(25) 
                           => n_1059, address_to_dram(24) => n_1060, 
                           address_to_dram(23) => n_1061, address_to_dram(22) 
                           => n_1062, address_to_dram(21) => n_1063, 
                           address_to_dram(20) => n_1064, address_to_dram(19) 
                           => n_1065, address_to_dram(18) => n_1066, 
                           address_to_dram(17) => n_1067, address_to_dram(16) 
                           => n_1068, address_to_dram(15) => n_1069, 
                           address_to_dram(14) => n_1070, address_to_dram(13) 
                           => n_1071, address_to_dram(12) => n_1072, 
                           address_to_dram(11) => n_1073, address_to_dram(10) 
                           => n_1074, address_to_dram(9) => n_1075, 
                           address_to_dram(8) => n_1076, address_to_dram(7) => 
                           n_1077, address_to_dram(6) => n_1078, 
                           address_to_dram(5) => n_1079, address_to_dram(4) => 
                           n_1080, address_to_dram(3) => n_1081, 
                           address_to_dram(2) => n_1082, address_to_dram(1) => 
                           n_1083, address_to_dram(0) => n_1084, 
                           data_to_dram(31) => n_1085, data_to_dram(30) => 
                           n_1086, data_to_dram(29) => n_1087, data_to_dram(28)
                           => n_1088, data_to_dram(27) => n_1089, 
                           data_to_dram(26) => n_1090, data_to_dram(25) => 
                           n_1091, data_to_dram(24) => n_1092, data_to_dram(23)
                           => n_1093, data_to_dram(22) => n_1094, 
                           data_to_dram(21) => n_1095, data_to_dram(20) => 
                           n_1096, data_to_dram(19) => n_1097, data_to_dram(18)
                           => n_1098, data_to_dram(17) => n_1099, 
                           data_to_dram(16) => n_1100, data_to_dram(15) => 
                           n_1101, data_to_dram(14) => n_1102, data_to_dram(13)
                           => n_1103, data_to_dram(12) => n_1104, 
                           data_to_dram(11) => n_1105, data_to_dram(10) => 
                           n_1106, data_to_dram(9) => n_1107, data_to_dram(8) 
                           => n_1108, data_to_dram(7) => n_1109, 
                           data_to_dram(6) => n_1110, data_to_dram(5) => n_1111
                           , data_to_dram(4) => n_1112, data_to_dram(3) => 
                           n_1113, data_to_dram(2) => n_1114, data_to_dram(1) 
                           => n_1115, data_to_dram(0) => n_1116, 
                           dram_to_dlx(31) => X_Logic0_port, dram_to_dlx(30) =>
                           X_Logic0_port, dram_to_dlx(29) => X_Logic0_port, 
                           dram_to_dlx(28) => X_Logic0_port, dram_to_dlx(27) =>
                           X_Logic0_port, dram_to_dlx(26) => X_Logic0_port, 
                           dram_to_dlx(25) => X_Logic0_port, dram_to_dlx(24) =>
                           X_Logic0_port, dram_to_dlx(23) => X_Logic0_port, 
                           dram_to_dlx(22) => X_Logic0_port, dram_to_dlx(21) =>
                           X_Logic0_port, dram_to_dlx(20) => X_Logic0_port, 
                           dram_to_dlx(19) => X_Logic0_port, dram_to_dlx(18) =>
                           X_Logic0_port, dram_to_dlx(17) => X_Logic0_port, 
                           dram_to_dlx(16) => X_Logic0_port, dram_to_dlx(15) =>
                           X_Logic0_port, dram_to_dlx(14) => X_Logic0_port, 
                           dram_to_dlx(13) => X_Logic0_port, dram_to_dlx(12) =>
                           X_Logic0_port, dram_to_dlx(11) => X_Logic0_port, 
                           dram_to_dlx(10) => X_Logic0_port, dram_to_dlx(9) => 
                           X_Logic0_port, dram_to_dlx(8) => X_Logic0_port, 
                           dram_to_dlx(7) => X_Logic0_port, dram_to_dlx(6) => 
                           X_Logic0_port, dram_to_dlx(5) => X_Logic0_port, 
                           dram_to_dlx(4) => X_Logic0_port, dram_to_dlx(3) => 
                           X_Logic0_port, dram_to_dlx(2) => X_Logic0_port, 
                           dram_to_dlx(1) => X_Logic0_port, dram_to_dlx(0) => 
                           X_Logic0_port, dram_we => n_1117, StallF => 
                           StallF_DP, StallD => StallD_DP, ForwardAD => 
                           ForwardAD_DP, ForwardBD => ForwardBD_DP, FlushE => 
                           FlushE_DP, rst_RF => rst, en_RF => X_Logic1_port, 
                           RsD_H(4) => RsD_H_DP_4_port, RsD_H(3) => 
                           RsD_H_DP_3_port, RsD_H(2) => RsD_H_DP_2_port, 
                           RsD_H(1) => RsD_H_DP_1_port, RsD_H(0) => 
                           RsD_H_DP_0_port, RtD_H(4) => RtD_H_DP_4_port, 
                           RtD_H(3) => RtD_H_DP_3_port, RtD_H(2) => 
                           RtD_H_DP_2_port, RtD_H(1) => RtD_H_DP_1_port, 
                           RtD_H(0) => RtD_H_DP_0_port, ForwardAE(1) => 
                           ForwardAE_DP_1_port, ForwardAE(0) => 
                           ForwardAE_DP_0_port, ForwardBE(1) => 
                           ForwardBE_DP_1_port, ForwardBE(0) => 
                           ForwardBE_DP_0_port, WriteRegE_H(4) => 
                           WriteRegE_H_DP_4_port, WriteRegE_H(3) => 
                           WriteRegE_H_DP_3_port, WriteRegE_H(2) => 
                           WriteRegE_H_DP_2_port, WriteRegE_H(1) => 
                           WriteRegE_H_DP_1_port, WriteRegE_H(0) => 
                           WriteRegE_H_DP_0_port, RsE_H(4) => RsE_H_DP_4_port, 
                           RsE_H(3) => RsE_H_DP_3_port, RsE_H(2) => 
                           RsE_H_DP_2_port, RsE_H(1) => RsE_H_DP_1_port, 
                           RsE_H(0) => RsE_H_DP_0_port, RtE_H(4) => 
                           RtE_H_DP_4_port, RtE_H(3) => RtE_H_DP_3_port, 
                           RtE_H(2) => RtE_H_DP_2_port, RtE_H(1) => 
                           RtE_H_DP_1_port, RtE_H(0) => RtE_H_DP_0_port, 
                           WriteRegMOut_H(4) => WriteRegMOut_H_DP_4_port, 
                           WriteRegMOut_H(3) => WriteRegMOut_H_DP_3_port, 
                           WriteRegMOut_H(2) => WriteRegMOut_H_DP_2_port, 
                           WriteRegMOut_H(1) => WriteRegMOut_H_DP_1_port, 
                           WriteRegMOut_H(0) => WriteRegMOut_H_DP_0_port, 
                           rst_mem => rst, WriteRegWBOut_H(4) => 
                           WriteRegWBOut_H_DP_4_port, WriteRegWBOut_H(3) => 
                           WriteRegWBOut_H_DP_3_port, WriteRegWBOut_H(2) => 
                           WriteRegWBOut_H_DP_2_port, WriteRegWBOut_H(1) => 
                           WriteRegWBOut_H_DP_1_port, WriteRegWBOut_H(0) => 
                           WriteRegWBOut_H_DP_0_port, OP(5) => OP_DP_5_port, 
                           OP(4) => OP_DP_4_port, OP(3) => OP_DP_3_port, OP(2) 
                           => OP_DP_2_port, OP(1) => OP_DP_1_port, OP(0) => 
                           OP_DP_0_port, FUNC(10) => FUNC_DP_10_port, FUNC(9) 
                           => FUNC_DP_9_port, FUNC(8) => FUNC_DP_8_port, 
                           FUNC(7) => FUNC_DP_7_port, FUNC(6) => FUNC_DP_6_port
                           , FUNC(5) => FUNC_DP_5_port, FUNC(4) => 
                           FUNC_DP_4_port, FUNC(3) => FUNC_DP_3_port, FUNC(2) 
                           => FUNC_DP_2_port, FUNC(1) => FUNC_DP_1_port, 
                           FUNC(0) => FUNC_DP_0_port, EqualD => EqualD_DP, FILL
                           => n_1118, SPILL => n_1119, PCSrcD => n2, RegWriteW 
                           => RegWriteW_CU, Select_ext => n2, CALL => n2, RET 
                           => n2, RD1_EN => n2, RD2_EN => n2, isJal => n2, 
                           Comp_control(1) => n2, Comp_control(0) => n2, 
                           RegDstE => n1, ALUSrcE => n1, ALUControlE(5) => n1, 
                           ALUControlE(4) => n1, ALUControlE(3) => n1, 
                           ALUControlE(2) => n1, ALUControlE(1) => n1, 
                           ALUControlE(0) => n1, en_ALU => n1, MemWriteM => 
                           MemWriteM_CU, MemToRegW => MemToRegW_CU);
   HazardUnit : hazard_detection_unit port map( RsD(4) => RsD_H_DP_4_port, 
                           RsD(3) => RsD_H_DP_3_port, RsD(2) => RsD_H_DP_2_port
                           , RsD(1) => RsD_H_DP_1_port, RsD(0) => 
                           RsD_H_DP_0_port, RtD(4) => RtD_H_DP_4_port, RtD(3) 
                           => RtD_H_DP_3_port, RtD(2) => RtD_H_DP_2_port, 
                           RtD(1) => RtD_H_DP_1_port, RtD(0) => RtD_H_DP_0_port
                           , RsE(4) => RsE_H_DP_4_port, RsE(3) => 
                           RsE_H_DP_3_port, RsE(2) => RsE_H_DP_2_port, RsE(1) 
                           => RsE_H_DP_1_port, RsE(0) => RsE_H_DP_0_port, 
                           RtE(4) => RtE_H_DP_4_port, RtE(3) => RtE_H_DP_3_port
                           , RtE(2) => RtE_H_DP_2_port, RtE(1) => 
                           RtE_H_DP_1_port, RtE(0) => RtE_H_DP_0_port, 
                           WriteRegM(4) => WriteRegMOut_H_DP_4_port, 
                           WriteRegM(3) => WriteRegMOut_H_DP_3_port, 
                           WriteRegM(2) => WriteRegMOut_H_DP_2_port, 
                           WriteRegM(1) => WriteRegMOut_H_DP_1_port, 
                           WriteRegM(0) => WriteRegMOut_H_DP_0_port, 
                           WriteRegW(4) => WriteRegWBOut_H_DP_4_port, 
                           WriteRegW(3) => WriteRegWBOut_H_DP_3_port, 
                           WriteRegW(2) => WriteRegWBOut_H_DP_2_port, 
                           WriteRegW(1) => WriteRegWBOut_H_DP_1_port, 
                           WriteRegW(0) => WriteRegWBOut_H_DP_0_port, 
                           WriteRegE(4) => WriteRegE_H_DP_4_port, WriteRegE(3) 
                           => WriteRegE_H_DP_3_port, WriteRegE(2) => 
                           WriteRegE_H_DP_2_port, WriteRegE(1) => 
                           WriteRegE_H_DP_1_port, WriteRegE(0) => 
                           WriteRegE_H_DP_0_port, BranchD => n2, MemToRegE => 
                           n1, MemToRegM => MemToRegM_H_CU, RegWriteM => 
                           RegWriteM_H_CU, RegWriteW => RegWriteW_H_CU, 
                           RegWriteE => n1, ForwardAD => ForwardAD_DP, 
                           ForwardBD => ForwardBD_DP, ForwardAE(1) => 
                           ForwardAE_DP_1_port, ForwardAE(0) => 
                           ForwardAE_DP_0_port, ForwardBE(1) => 
                           ForwardBE_DP_1_port, ForwardBE(0) => 
                           ForwardBE_DP_0_port, StallF => StallF_DP, StallD => 
                           StallD_DP, FlushE => n_1120);
   n1 <= '0';
   n2 <= '0';
   FlushE_DP <= '0';

end SYN_Behavioral;
